//
// Verilog description for cell lab_7_top, 
// 07/07/23 00:04:51
//
// Precision RTL Synthesis, 64-bit 2018.1.0.19//


module lab_7_top ( clk, reset, key_in, data_in, load, data_out ) ;

    input clk ;
    input reset ;
    input [63:0]key_in ;
    input [63:0]data_in ;
    input load ;
    output [63:0]data_out ;

    wire [63:0]data_out_1_0;
    wire \plaintext(63)  , \plaintext(39)  , \plaintext(37)  , \plaintext(5)  , 
         \key_samp(63)  , \key_samp(62)  , \key_samp(61)  , \key_samp(60)  , 
         \key_samp(59)  , \key_samp(58)  , \key_samp(57)  , \key_samp(55)  , 
         \key_samp(54)  , \key_samp(53)  , \key_samp(52)  , \key_samp(51)  , 
         \key_samp(50)  , \key_samp(49)  , \key_samp(47)  , \key_samp(46)  , 
         \key_samp(45)  , \key_samp(44)  , \key_samp(43)  , \key_samp(42)  , 
         \key_samp(41)  , \key_samp(39)  , \key_samp(38)  , \key_samp(37)  , 
         \key_samp(36)  , \key_samp(35)  , \key_samp(34)  , \key_samp(33)  , 
         \key_samp(31)  , \key_samp(30)  , \key_samp(29)  , \key_samp(28)  , 
         \key_samp(27)  , \key_samp(26)  , \key_samp(25)  , \key_samp(23)  , 
         \key_samp(22)  , \key_samp(21)  , \key_samp(20)  , \key_samp(19)  , 
         \key_samp(18)  , \key_samp(17)  , \key_samp(15)  , \key_samp(14)  , 
         \key_samp(13)  , \key_samp(12)  , \key_samp(11)  , \key_samp(10)  , 
         \key_samp(9)  , \key_samp(7)  , \key_samp(6)  , \key_samp(5)  , 
         \key_samp(4)  , \key_samp(3)  , \key_samp(2)  , \key_samp(1)  ;
    wire clk_int;
    wire reset_int;
    wire [63:8]key_in_int;
    wire [63:0]data_in_int;
    wire load_int, nx7754z1, nx5760z1, nx3766z1, nx1772z1, nx65314z1, nx55009z1, 
         nx53015z1, nx51021z1, nx49027z1, nx47033z1, nx44040z1, nx42046z1, 
         nx40052z1, nx38058z1, nx36064z1, nx33071z1, nx31077z1, nx29083z1, 
         nx27089z1, nx25095z1, nx22102z1, nx20108z1, nx18114z1, nx16120z1, 
         nx14126z1, nx11133z1, nx9139z1, nx7145z1, nx5151z1, nx3157z1, nx164z1, 
         nx63706z1, nx41410z1, nx61354z1, nx21466z1, nx45398z1, nx63348z1, 
         nx50385z1, nx34429z1, nx65342z1, nx23460z1, nx26453z1, nx39416z1, 
         nx37422z1, nx28447z1, nx22549z1, nx52379z1, nx6787z1, nx16567z1, 
         nx17478z1, nx32435z1, nx14573z1, nx54373z1, nx48391z1, nx4793z1, 
         nx1800z1, nx15484z1, nx19472z1, nx30441z1, nx43404z1, nx56367z1, 
         nx59360z1, nx20555z1, nx18561z1, nx15286z132, nx5589z279, nx15286z131, 
         nx5589z274, nx15286z130, nx5589z269, nx15286z160, nx15286z159, 
         nx15286z158, nx15286z157, nx15286z163, nx15286z162, nx15286z161, 
         nx15286z164, nx15286z153, nx5589z249, nx15286z154, nx5589z259, 
         nx15286z155, nx15286z156, nx15286z144, nx15286z143, nx15286z142, 
         nx15286z141, nx15286z145, nx5589z234, nx15286z146, nx5589z239, 
         nx15286z147, nx15286z148, nx15286z133, nx5589z224, nx15286z135, 
         nx5589z219, nx15286z134, nx5589z199, nx15286z136, nx5589z214, 
         nx15286z149, nx5589z229, nx15286z126, nx15286z127, nx15286z128, 
         nx15286z129, nx15286z150, nx5589z254, nx15286z151, nx5589z264, 
         nx15286z152, nx15286z110, nx15286z111, nx15286z112, nx15286z113, 
         nx15286z137, nx5589z209, nx15286z118, nx5589z280, nx15286z119, 
         nx15286z120, nx15286z121, nx5589z182, nx15286z138, nx5589z189, 
         nx15286z106, nx15286z107, nx15286z108, nx5589z275, nx15286z109, 
         nx5589z145, nx15286z114, nx5589z177, nx15286z115, nx5589z172, 
         nx15286z116, nx5589z152, nx15286z117, nx5589z167, nx15286z122, 
         nx15286z124, nx15286z123, nx5589z138, nx15286z125, nx5589z270, 
         nx15286z139, nx5589z204, nx15286z98, nx5589z162, nx15286z99, 
         nx15286z100, nx15286z101, nx5589z157, nx15286z87, nx15286z88, 
         nx15286z89, nx15286z140, nx5589z194, nx5589z244, nx15286z104, 
         nx5589z128, nx15286z94, nx15286z95, nx15286z103, nx5589z133, nx15286z92, 
         nx5589z250, nx15286z93, nx5589z260, nx15286z105, nx5589z118, nx15286z90, 
         nx5589z235, nx15286z91, nx5589z240, nx5589z255, nx5589z230, nx15286z97, 
         nx5589z265, nx15286z70, nx15286z69, nx15286z96, nx15286z102, nx5589z123, 
         nx5589z220, nx5589z225, nx5589z215, nx15286z74, nx15286z75, nx15286z76, 
         nx5589z200, nx5589z205, nx15286z64, nx15286z65, nx5589z163, nx15286z66, 
         nx15286z67, nx5589z158, nx15286z84, nx5589z210, nx15286z81, nx5589z183, 
         nx15286z82, nx5589z281, nx15286z83, nx5589z178, nx5589z168, nx15286z79, 
         nx5589z173, nx15286z80, nx5589z153, nx15286z86, nx5589z190, nx5589z146, 
         nx15286z68, nx5589z276, nx15286z77, nx15286z44, nx15286z45, nx15286z46, 
         nx15286z47, nx5589z139, nx5589z271, nx15286z42, nx15286z41, nx15286z43, 
         nx15286z40, nx15286z78, nx15286z85, nx5589z195, nx5589z245, nx15286z72, 
         nx5589z129, nx15286z48, nx15286z49, nx15286z50, nx15286z51, nx5589z119, 
         nx15286z60, nx5589z236, nx15286z61, nx15286z62, nx15286z63, nx5589z241, 
         nx15286z71, nx5589z134, nx15286z56, nx5589z251, nx15286z57, nx15286z58, 
         nx15286z59, nx5589z261, nx15286z54, nx5589z256, nx15286z53, nx5589z266, 
         nx15286z52, nx15286z55, nx5589z231, nx15286z14, nx15286z16, nx15286z15, 
         nx15286z73, nx5589z124, nx15286z32, nx5589z216, nx15286z17, nx15286z18, 
         nx15286z19, nx15286z20, nx15286z35, nx5589z221, nx15286z34, nx5589z226, 
         nx15286z33, nx5589z201, nx15286z36, nx5589z191, nx15286z6, nx15286z7, 
         nx15286z24, nx5589z174, nx15286z25, nx5589z179, nx15286z26, nx5589z169, 
         nx15286z27, nx5589z154, nx15286z37, nx5589z206, nx15286z8, nx5589z164, 
         nx15286z9, nx5589z159, nx15286z10, nx15286z21, nx5589z272, nx5589z273, 
         nx15286z22, nx5589z140, nx15286z23, nx15286z38, nx5589z211, nx15286z28, 
         nx5589z184, nx15286z29, nx5589z277, nx5589z278, nx15286z30, nx5589z282, 
         nx5589z283, nx15286z31, nx5589z147, nx15286z39, nx5589z196, nx5589z246, 
         nx15286z12, nx5589z135, nx5589z262, nx5589z263, nx5589z252, nx5589z253, 
         nx15286z13, nx5589z130, nx15286z11, nx5589z120, nx5589z242, nx5589z243, 
         nx5589z237, nx5589z238, nx5589z257, nx5589z258, nx5589z267, nx5589z268, 
         nx5589z232, nx5589z233, nx5589z125, nx5589z217, nx5589z218, nx5589z222, 
         nx5589z223, nx5589z227, nx5589z228, nx5589z202, nx5589z203, nx5589z212, 
         nx5589z185, nx5589z186, nx5589z187, nx5589z188, nx5589z213, nx5589z192, 
         nx5589z150, nx5589z151, nx5589z148, nx5589z149, nx5589z193, nx5589z143, 
         nx5589z144, nx5589z141, nx5589z142, nx5589z197, nx5589z198, nx5589z175, 
         nx5589z176, nx5589z180, nx5589z181, nx5589z170, nx5589z171, nx5589z155, 
         nx5589z156, nx5589z207, nx5589z165, nx5589z166, nx5589z160, nx5589z161, 
         nx5589z208, nx5589z247, nx5589z131, nx5589z132, nx5589z136, nx5589z104, 
         nx5589z105, nx5589z116, nx5589z117, nx5589z137, nx5589z121, nx5589z100, 
         nx5589z101, nx5589z102, nx5589z103, nx5589z122, nx5589z126, nx5589z106, 
         nx5589z107, nx5589z36, nx5589z43, nx5589z110, nx5589z111, nx5589z127, 
         nx5589z114, nx5589z115, nx5589z69, nx5589z112, nx5589z113, nx5589z76, 
         nx5589z77, nx5589z53, nx5589z54, nx5589z46, nx5589z98, nx5589z99, 
         nx5589z82, nx5589z83, nx5589z108, nx5589z92, nx5589z93, nx5589z78, 
         nx5589z79, nx5589z88, nx5589z89, nx5589z80, nx5589z81, nx5589z109, 
         nx5589z19, nx5589z96, nx5589z97, nx5589z90, nx5589z91, nx5589z11, 
         nx5589z16, nx5589z248, nx5589z94, nx5589z84, nx5589z67, nx5589z68, 
         nx5589z65, nx5589z66, nx5589z85, nx5589z55, nx5589z56, nx5589z86, 
         nx5589z51, nx5589z52, nx5589z44, nx5589z45, nx5589z87, nx5589z61, 
         nx5589z62, nx5589z63, nx5589z64, nx5589z70, nx5589z71, nx5589z74, 
         nx5589z34, nx5589z35, nx5589z59, nx5589z60, nx5589z37, nx5589z38, 
         nx5589z57, nx5589z58, nx5589z75, nx5589z49, nx5589z26, nx5589z27, 
         nx5589z24, nx5589z25, nx5589z50, nx5589z41, nx5589z3, nx5589z4, 
         nx5589z14, nx5589z15, nx5589z42, nx5589z39, nx5589z40, nx5589z47, 
         nx5589z30, nx5589z31, nx5589z32, nx5589z33, nx5589z48, nx5589z17, 
         nx5589z18, nx5589z20, nx5589z21, nx15286z4, nx5589z28, nx5589z29, 
         nx5589z12, nx5589z13, nx5589z22, nx5589z23, nx5589z95, nx5589z72, 
         nx5589z7, nx5589z8, nx5589z9, nx15286z5, nx5589z1, nx5589z10, nx5589z5, 
         nx5589z6, nx5589z2, nx15286z1, nx15286z2, nx5589z73, nx15286z3, nx4;



    OBUF \data_out_obuf(0)  (.O (data_out[0]), .I (data_out_1_0[0])) ;
    OBUF \data_out_obuf(1)  (.O (data_out[1]), .I (data_out_1_0[1])) ;
    OBUF \data_out_obuf(2)  (.O (data_out[2]), .I (data_out_1_0[2])) ;
    OBUF \data_out_obuf(3)  (.O (data_out[3]), .I (data_out_1_0[3])) ;
    OBUF \data_out_obuf(4)  (.O (data_out[4]), .I (data_out_1_0[4])) ;
    OBUF \data_out_obuf(5)  (.O (data_out[5]), .I (data_out_1_0[5])) ;
    OBUF \data_out_obuf(6)  (.O (data_out[6]), .I (data_out_1_0[6])) ;
    OBUF \data_out_obuf(7)  (.O (data_out[7]), .I (data_out_1_0[7])) ;
    OBUF \data_out_obuf(8)  (.O (data_out[8]), .I (data_out_1_0[8])) ;
    OBUF \data_out_obuf(9)  (.O (data_out[9]), .I (data_out_1_0[9])) ;
    OBUF \data_out_obuf(10)  (.O (data_out[10]), .I (data_out_1_0[10])) ;
    OBUF \data_out_obuf(11)  (.O (data_out[11]), .I (data_out_1_0[11])) ;
    OBUF \data_out_obuf(12)  (.O (data_out[12]), .I (data_out_1_0[12])) ;
    OBUF \data_out_obuf(13)  (.O (data_out[13]), .I (data_out_1_0[13])) ;
    OBUF \data_out_obuf(14)  (.O (data_out[14]), .I (data_out_1_0[14])) ;
    OBUF \data_out_obuf(15)  (.O (data_out[15]), .I (data_out_1_0[15])) ;
    OBUF \data_out_obuf(16)  (.O (data_out[16]), .I (data_out_1_0[16])) ;
    OBUF \data_out_obuf(17)  (.O (data_out[17]), .I (data_out_1_0[17])) ;
    OBUF \data_out_obuf(18)  (.O (data_out[18]), .I (data_out_1_0[18])) ;
    OBUF \data_out_obuf(19)  (.O (data_out[19]), .I (data_out_1_0[19])) ;
    OBUF \data_out_obuf(20)  (.O (data_out[20]), .I (data_out_1_0[20])) ;
    OBUF \data_out_obuf(21)  (.O (data_out[21]), .I (data_out_1_0[21])) ;
    OBUF \data_out_obuf(22)  (.O (data_out[22]), .I (data_out_1_0[22])) ;
    OBUF \data_out_obuf(23)  (.O (data_out[23]), .I (data_out_1_0[23])) ;
    OBUF \data_out_obuf(24)  (.O (data_out[24]), .I (data_out_1_0[24])) ;
    OBUF \data_out_obuf(25)  (.O (data_out[25]), .I (data_out_1_0[25])) ;
    OBUF \data_out_obuf(26)  (.O (data_out[26]), .I (data_out_1_0[26])) ;
    OBUF \data_out_obuf(27)  (.O (data_out[27]), .I (data_out_1_0[27])) ;
    OBUF \data_out_obuf(28)  (.O (data_out[28]), .I (data_out_1_0[28])) ;
    OBUF \data_out_obuf(29)  (.O (data_out[29]), .I (data_out_1_0[29])) ;
    OBUF \data_out_obuf(30)  (.O (data_out[30]), .I (data_out_1_0[30])) ;
    OBUF \data_out_obuf(31)  (.O (data_out[31]), .I (data_out_1_0[31])) ;
    OBUF \data_out_obuf(32)  (.O (data_out[32]), .I (data_out_1_0[32])) ;
    OBUF \data_out_obuf(33)  (.O (data_out[33]), .I (data_out_1_0[33])) ;
    OBUF \data_out_obuf(34)  (.O (data_out[34]), .I (data_out_1_0[34])) ;
    OBUF \data_out_obuf(35)  (.O (data_out[35]), .I (data_out_1_0[35])) ;
    OBUF \data_out_obuf(36)  (.O (data_out[36]), .I (data_out_1_0[36])) ;
    OBUF \data_out_obuf(37)  (.O (data_out[37]), .I (data_out_1_0[37])) ;
    OBUF \data_out_obuf(38)  (.O (data_out[38]), .I (data_out_1_0[38])) ;
    OBUF \data_out_obuf(39)  (.O (data_out[39]), .I (data_out_1_0[39])) ;
    OBUF \data_out_obuf(40)  (.O (data_out[40]), .I (data_out_1_0[40])) ;
    OBUF \data_out_obuf(41)  (.O (data_out[41]), .I (data_out_1_0[41])) ;
    OBUF \data_out_obuf(42)  (.O (data_out[42]), .I (data_out_1_0[42])) ;
    OBUF \data_out_obuf(43)  (.O (data_out[43]), .I (data_out_1_0[43])) ;
    OBUF \data_out_obuf(44)  (.O (data_out[44]), .I (data_out_1_0[44])) ;
    OBUF \data_out_obuf(45)  (.O (data_out[45]), .I (data_out_1_0[45])) ;
    OBUF \data_out_obuf(46)  (.O (data_out[46]), .I (data_out_1_0[46])) ;
    OBUF \data_out_obuf(47)  (.O (data_out[47]), .I (data_out_1_0[47])) ;
    OBUF \data_out_obuf(48)  (.O (data_out[48]), .I (data_out_1_0[48])) ;
    OBUF \data_out_obuf(49)  (.O (data_out[49]), .I (data_out_1_0[49])) ;
    OBUF \data_out_obuf(50)  (.O (data_out[50]), .I (data_out_1_0[50])) ;
    OBUF \data_out_obuf(51)  (.O (data_out[51]), .I (data_out_1_0[51])) ;
    OBUF \data_out_obuf(52)  (.O (data_out[52]), .I (data_out_1_0[52])) ;
    OBUF \data_out_obuf(53)  (.O (data_out[53]), .I (data_out_1_0[53])) ;
    OBUF \data_out_obuf(54)  (.O (data_out[54]), .I (data_out_1_0[54])) ;
    OBUF \data_out_obuf(55)  (.O (data_out[55]), .I (data_out_1_0[55])) ;
    OBUF \data_out_obuf(56)  (.O (data_out[56]), .I (data_out_1_0[56])) ;
    OBUF \data_out_obuf(57)  (.O (data_out[57]), .I (data_out_1_0[57])) ;
    OBUF \data_out_obuf(58)  (.O (data_out[58]), .I (data_out_1_0[58])) ;
    OBUF \data_out_obuf(59)  (.O (data_out[59]), .I (data_out_1_0[59])) ;
    OBUF \data_out_obuf(60)  (.O (data_out[60]), .I (data_out_1_0[60])) ;
    OBUF \data_out_obuf(61)  (.O (data_out[61]), .I (data_out_1_0[61])) ;
    OBUF \data_out_obuf(62)  (.O (data_out[62]), .I (data_out_1_0[62])) ;
    OBUF \data_out_obuf(63)  (.O (data_out[63]), .I (data_out_1_0[63])) ;
    IBUF load_ibuf (.O (load_int), .I (load)) ;
    IBUF \data_in_ibuf(0)  (.O (data_in_int[0]), .I (data_in[0])) ;
    IBUF \data_in_ibuf(1)  (.O (data_in_int[1]), .I (data_in[1])) ;
    IBUF \data_in_ibuf(2)  (.O (data_in_int[2]), .I (data_in[2])) ;
    IBUF \data_in_ibuf(3)  (.O (data_in_int[3]), .I (data_in[3])) ;
    IBUF \data_in_ibuf(4)  (.O (data_in_int[4]), .I (data_in[4])) ;
    IBUF \data_in_ibuf(5)  (.O (data_in_int[5]), .I (data_in[5])) ;
    IBUF \data_in_ibuf(6)  (.O (data_in_int[6]), .I (data_in[6])) ;
    IBUF \data_in_ibuf(7)  (.O (data_in_int[7]), .I (data_in[7])) ;
    IBUF \data_in_ibuf(8)  (.O (data_in_int[8]), .I (data_in[8])) ;
    IBUF \data_in_ibuf(9)  (.O (data_in_int[9]), .I (data_in[9])) ;
    IBUF \data_in_ibuf(10)  (.O (data_in_int[10]), .I (data_in[10])) ;
    IBUF \data_in_ibuf(11)  (.O (data_in_int[11]), .I (data_in[11])) ;
    IBUF \data_in_ibuf(12)  (.O (data_in_int[12]), .I (data_in[12])) ;
    IBUF \data_in_ibuf(13)  (.O (data_in_int[13]), .I (data_in[13])) ;
    IBUF \data_in_ibuf(14)  (.O (data_in_int[14]), .I (data_in[14])) ;
    IBUF \data_in_ibuf(15)  (.O (data_in_int[15]), .I (data_in[15])) ;
    IBUF \data_in_ibuf(16)  (.O (data_in_int[16]), .I (data_in[16])) ;
    IBUF \data_in_ibuf(17)  (.O (data_in_int[17]), .I (data_in[17])) ;
    IBUF \data_in_ibuf(18)  (.O (data_in_int[18]), .I (data_in[18])) ;
    IBUF \data_in_ibuf(19)  (.O (data_in_int[19]), .I (data_in[19])) ;
    IBUF \data_in_ibuf(20)  (.O (data_in_int[20]), .I (data_in[20])) ;
    IBUF \data_in_ibuf(21)  (.O (data_in_int[21]), .I (data_in[21])) ;
    IBUF \data_in_ibuf(22)  (.O (data_in_int[22]), .I (data_in[22])) ;
    IBUF \data_in_ibuf(23)  (.O (data_in_int[23]), .I (data_in[23])) ;
    IBUF \data_in_ibuf(24)  (.O (data_in_int[24]), .I (data_in[24])) ;
    IBUF \data_in_ibuf(25)  (.O (data_in_int[25]), .I (data_in[25])) ;
    IBUF \data_in_ibuf(26)  (.O (data_in_int[26]), .I (data_in[26])) ;
    IBUF \data_in_ibuf(27)  (.O (data_in_int[27]), .I (data_in[27])) ;
    IBUF \data_in_ibuf(28)  (.O (data_in_int[28]), .I (data_in[28])) ;
    IBUF \data_in_ibuf(29)  (.O (data_in_int[29]), .I (data_in[29])) ;
    IBUF \data_in_ibuf(30)  (.O (data_in_int[30]), .I (data_in[30])) ;
    IBUF \data_in_ibuf(31)  (.O (data_in_int[31]), .I (data_in[31])) ;
    IBUF \data_in_ibuf(32)  (.O (data_in_int[32]), .I (data_in[32])) ;
    IBUF \data_in_ibuf(33)  (.O (data_in_int[33]), .I (data_in[33])) ;
    IBUF \data_in_ibuf(34)  (.O (data_in_int[34]), .I (data_in[34])) ;
    IBUF \data_in_ibuf(35)  (.O (data_in_int[35]), .I (data_in[35])) ;
    IBUF \data_in_ibuf(36)  (.O (data_in_int[36]), .I (data_in[36])) ;
    IBUF \data_in_ibuf(37)  (.O (data_in_int[37]), .I (data_in[37])) ;
    IBUF \data_in_ibuf(38)  (.O (data_in_int[38]), .I (data_in[38])) ;
    IBUF \data_in_ibuf(39)  (.O (data_in_int[39]), .I (data_in[39])) ;
    IBUF \data_in_ibuf(40)  (.O (data_in_int[40]), .I (data_in[40])) ;
    IBUF \data_in_ibuf(41)  (.O (data_in_int[41]), .I (data_in[41])) ;
    IBUF \data_in_ibuf(42)  (.O (data_in_int[42]), .I (data_in[42])) ;
    IBUF \data_in_ibuf(43)  (.O (data_in_int[43]), .I (data_in[43])) ;
    IBUF \data_in_ibuf(44)  (.O (data_in_int[44]), .I (data_in[44])) ;
    IBUF \data_in_ibuf(45)  (.O (data_in_int[45]), .I (data_in[45])) ;
    IBUF \data_in_ibuf(46)  (.O (data_in_int[46]), .I (data_in[46])) ;
    IBUF \data_in_ibuf(47)  (.O (data_in_int[47]), .I (data_in[47])) ;
    IBUF \data_in_ibuf(48)  (.O (data_in_int[48]), .I (data_in[48])) ;
    IBUF \data_in_ibuf(49)  (.O (data_in_int[49]), .I (data_in[49])) ;
    IBUF \data_in_ibuf(50)  (.O (data_in_int[50]), .I (data_in[50])) ;
    IBUF \data_in_ibuf(51)  (.O (data_in_int[51]), .I (data_in[51])) ;
    IBUF \data_in_ibuf(52)  (.O (data_in_int[52]), .I (data_in[52])) ;
    IBUF \data_in_ibuf(53)  (.O (data_in_int[53]), .I (data_in[53])) ;
    IBUF \data_in_ibuf(54)  (.O (data_in_int[54]), .I (data_in[54])) ;
    IBUF \data_in_ibuf(55)  (.O (data_in_int[55]), .I (data_in[55])) ;
    IBUF \data_in_ibuf(56)  (.O (data_in_int[56]), .I (data_in[56])) ;
    IBUF \data_in_ibuf(57)  (.O (data_in_int[57]), .I (data_in[57])) ;
    IBUF \data_in_ibuf(58)  (.O (data_in_int[58]), .I (data_in[58])) ;
    IBUF \data_in_ibuf(59)  (.O (data_in_int[59]), .I (data_in[59])) ;
    IBUF \data_in_ibuf(60)  (.O (data_in_int[60]), .I (data_in[60])) ;
    IBUF \data_in_ibuf(61)  (.O (data_in_int[61]), .I (data_in[61])) ;
    IBUF \data_in_ibuf(62)  (.O (data_in_int[62]), .I (data_in[62])) ;
    IBUF \data_in_ibuf(63)  (.O (data_in_int[63]), .I (data_in[63])) ;
    IBUF \key_in_ibuf(1)  (.O (key_in_int[8]), .I (key_in[1])) ;
    IBUF \key_in_ibuf(2)  (.O (key_in_int[9]), .I (key_in[2])) ;
    IBUF \key_in_ibuf(3)  (.O (key_in_int[10]), .I (key_in[3])) ;
    IBUF \key_in_ibuf(4)  (.O (key_in_int[11]), .I (key_in[4])) ;
    IBUF \key_in_ibuf(5)  (.O (key_in_int[12]), .I (key_in[5])) ;
    IBUF \key_in_ibuf(6)  (.O (key_in_int[13]), .I (key_in[6])) ;
    IBUF \key_in_ibuf(7)  (.O (key_in_int[14]), .I (key_in[7])) ;
    IBUF \key_in_ibuf(9)  (.O (key_in_int[15]), .I (key_in[9])) ;
    IBUF \key_in_ibuf(10)  (.O (key_in_int[16]), .I (key_in[10])) ;
    IBUF \key_in_ibuf(11)  (.O (key_in_int[17]), .I (key_in[11])) ;
    IBUF \key_in_ibuf(12)  (.O (key_in_int[18]), .I (key_in[12])) ;
    IBUF \key_in_ibuf(13)  (.O (key_in_int[19]), .I (key_in[13])) ;
    IBUF \key_in_ibuf(14)  (.O (key_in_int[20]), .I (key_in[14])) ;
    IBUF \key_in_ibuf(15)  (.O (key_in_int[21]), .I (key_in[15])) ;
    IBUF \key_in_ibuf(17)  (.O (key_in_int[22]), .I (key_in[17])) ;
    IBUF \key_in_ibuf(18)  (.O (key_in_int[23]), .I (key_in[18])) ;
    IBUF \key_in_ibuf(19)  (.O (key_in_int[24]), .I (key_in[19])) ;
    IBUF \key_in_ibuf(20)  (.O (key_in_int[25]), .I (key_in[20])) ;
    IBUF \key_in_ibuf(21)  (.O (key_in_int[26]), .I (key_in[21])) ;
    IBUF \key_in_ibuf(22)  (.O (key_in_int[27]), .I (key_in[22])) ;
    IBUF \key_in_ibuf(23)  (.O (key_in_int[28]), .I (key_in[23])) ;
    IBUF \key_in_ibuf(25)  (.O (key_in_int[29]), .I (key_in[25])) ;
    IBUF \key_in_ibuf(26)  (.O (key_in_int[30]), .I (key_in[26])) ;
    IBUF \key_in_ibuf(27)  (.O (key_in_int[31]), .I (key_in[27])) ;
    IBUF \key_in_ibuf(28)  (.O (key_in_int[32]), .I (key_in[28])) ;
    IBUF \key_in_ibuf(29)  (.O (key_in_int[33]), .I (key_in[29])) ;
    IBUF \key_in_ibuf(30)  (.O (key_in_int[34]), .I (key_in[30])) ;
    IBUF \key_in_ibuf(31)  (.O (key_in_int[35]), .I (key_in[31])) ;
    IBUF \key_in_ibuf(33)  (.O (key_in_int[36]), .I (key_in[33])) ;
    IBUF \key_in_ibuf(34)  (.O (key_in_int[37]), .I (key_in[34])) ;
    IBUF \key_in_ibuf(35)  (.O (key_in_int[38]), .I (key_in[35])) ;
    IBUF \key_in_ibuf(36)  (.O (key_in_int[39]), .I (key_in[36])) ;
    IBUF \key_in_ibuf(37)  (.O (key_in_int[40]), .I (key_in[37])) ;
    IBUF \key_in_ibuf(38)  (.O (key_in_int[41]), .I (key_in[38])) ;
    IBUF \key_in_ibuf(39)  (.O (key_in_int[42]), .I (key_in[39])) ;
    IBUF \key_in_ibuf(41)  (.O (key_in_int[43]), .I (key_in[41])) ;
    IBUF \key_in_ibuf(42)  (.O (key_in_int[44]), .I (key_in[42])) ;
    IBUF \key_in_ibuf(43)  (.O (key_in_int[45]), .I (key_in[43])) ;
    IBUF \key_in_ibuf(44)  (.O (key_in_int[46]), .I (key_in[44])) ;
    IBUF \key_in_ibuf(45)  (.O (key_in_int[47]), .I (key_in[45])) ;
    IBUF \key_in_ibuf(46)  (.O (key_in_int[48]), .I (key_in[46])) ;
    IBUF \key_in_ibuf(47)  (.O (key_in_int[49]), .I (key_in[47])) ;
    IBUF \key_in_ibuf(49)  (.O (key_in_int[50]), .I (key_in[49])) ;
    IBUF \key_in_ibuf(50)  (.O (key_in_int[51]), .I (key_in[50])) ;
    IBUF \key_in_ibuf(51)  (.O (key_in_int[52]), .I (key_in[51])) ;
    IBUF \key_in_ibuf(52)  (.O (key_in_int[53]), .I (key_in[52])) ;
    IBUF \key_in_ibuf(53)  (.O (key_in_int[54]), .I (key_in[53])) ;
    IBUF \key_in_ibuf(54)  (.O (key_in_int[55]), .I (key_in[54])) ;
    IBUF \key_in_ibuf(55)  (.O (key_in_int[56]), .I (key_in[55])) ;
    IBUF \key_in_ibuf(57)  (.O (key_in_int[57]), .I (key_in[57])) ;
    IBUF \key_in_ibuf(58)  (.O (key_in_int[58]), .I (key_in[58])) ;
    IBUF \key_in_ibuf(59)  (.O (key_in_int[59]), .I (key_in[59])) ;
    IBUF \key_in_ibuf(60)  (.O (key_in_int[60]), .I (key_in[60])) ;
    IBUF \key_in_ibuf(61)  (.O (key_in_int[61]), .I (key_in[61])) ;
    IBUF \key_in_ibuf(62)  (.O (key_in_int[62]), .I (key_in[62])) ;
    IBUF \key_in_ibuf(63)  (.O (key_in_int[63]), .I (key_in[63])) ;
    IBUF reset_ibuf (.O (reset_int), .I (reset)) ;
    input_register_0 i_data_samp (.px3886 (nx5589z73), .px3870 (nx15286z1), .px3872 (
                     nx15286z2), .px3923 (nx15286z3), .px3761 (nx5589z6), .px3750 (
                     nx5589z10), .px3737 (nx5589z8), .px3717 (nx5589z23), .px3703 (
                     nx5589z29), .px3689 (nx5589z21), .px3675 (nx5589z18), .px3667 (
                     nx5589z48), .px3666 (nx5589z33), .px3658 (nx5589z31), .px3650 (
                     nx5589z40), .px3647 (nx5589z42), .px3639 (nx5589z15), .px3630 (
                     nx5589z50), .px3627 (nx5589z25), .px3697 (nx15286z4), .px3624 (
                     nx5589z27), .px3611 (nx5589z75), .px3607 (nx5589z58), .px3744 (
                     nx15286z5), .px3591 (nx5589z38), .px3588 (nx5589z60), .px3585 (
                     nx5589z35), .px3576 (nx5589z71), .px3563 (nx5589z64), .px3560 (
                     nx5589z62), .px3551 (nx5589z87), .px3547 (nx5589z45), .px3544 (
                     nx5589z52), .px3534 (nx5589z56), .px3515 (nx5589z66), .px3512 (
                     nx5589z68), .px3455 (nx5589z91), .px3452 (nx5589z97), .px3444 (
                     nx5589z109), .px3443 (nx5589z81), .px3434 (nx5589z93), .px3411 (
                     nx5589z99), .px3374 (nx5589z113), .px3739 (nx5589z9), .px3649 (
                     nx5589z39), .px3632 (nx5589z41), .px3523 (nx5589z55), .px3752 (
                     nx5589z5), .px3652 (nx5589z47), .px3546 (nx5589z44), .px3425 (
                     nx5589z108), .px3615 (nx5589z49), .px3543 (nx5589z51), .px3582 (
                     nx5589z74), .px3726 (nx5589z7), .px3584 (nx5589z34), .px3590 (
                     nx5589z37), .px3433 (nx5589z92), .px3626 (nx5589z24), .px3596 (
                     nx5589z57), .px3587 (nx5589z59), .px3559 (nx5589z61), .px3781 (
                     nx5589z2), .px3373 (nx5589z112), .px3562 (nx5589z63), .px3442 (
                     nx5589z80), .px3638 (nx5589z14), .px3623 (nx5589z26), .px3511 (
                     nx5589z67), .px3514 (nx5589z65), .px3745 (nx5589z1), .px3724 (
                     nx5589z72), .px3565 (nx5589z70), .px3674 (nx5589z17), .px3665 (
                     nx5589z32), .px3536 (nx5589z86), .px3410 (nx5589z98), .px3657 (
                     nx5589z30), .px3451 (nx5589z96), .px3702 (nx5589z28), .px3688 (
                     nx5589z20), .px3454 (nx5589z90), .px3716 (nx5589z22), .px3635 (
                     nx5589z3), .px3636 (nx5589z4), .px3705 (nx5589z12), .px3714 (
                     nx5589z13), .px2959 (nx15286z6), .px2963 (nx15286z7), .px2986 (
                     nx15286z8), .px2996 (nx15286z9), .px2999 (nx15286z10), .px3506 (
                     nx5589z84), .px3521 (nx5589z85), .px3089 (nx15286z11), .px3059 (
                     nx15286z12), .px3076 (nx15286z13), .px2921 (nx15286z14), .px2925 (
                     nx15286z15), .px2924 (nx15286z16), .px2933 (nx15286z17), .px2934 (
                     nx15286z18), .px2935 (nx15286z19), .px2939 (nx15286z20), .px3005 (
                     nx15286z21), .px3008 (nx15286z22), .px3015 (nx15286z23), .\p_key_samp(15)   (
                     \key_samp(15)  ), .px2966 (nx15286z24), .px2969 (nx15286z25
                     ), .px2972 (nx15286z26), .px2981 (nx15286z27), .px3021 (
                     nx15286z28), .px3034 (nx15286z29), .px3040 (nx15286z30), .px3053 (
                     nx15286z31), .px3436 (nx5589z78), .px3437 (nx5589z79), .px3483 (
                     nx5589z16), .px2928 (nx15286z32), .px2944 (nx15286z33), .px2942 (
                     nx15286z34), .px2940 (nx15286z35), .\p_key_samp(44)   (
                     \key_samp(44)  ), .px2952 (nx15286z36), .px2984 (nx15286z37
                     ), .px3016 (nx15286z38), .px3056 (nx15286z39), .px3439 (
                     nx5589z88), .px3440 (nx5589z89), .px2865 (nx15286z40), .px2859 (
                     nx15286z41), .px2858 (nx15286z42), .px2860 (nx15286z43), .px2844 (
                     nx15286z44), .px2845 (nx15286z45), .px2846 (nx15286z46), .px2847 (
                     nx15286z47), .\p_key_samp(50)   (\key_samp(50)  ), .px2872 (
                     nx15286z48), .px2877 (nx15286z49), .px2878 (nx15286z50), .px2879 (
                     nx15286z51), .px3448 (nx5589z19), .px2912 (nx15286z52), .px2908 (
                     nx15286z53), .px2906 (nx15286z54), .px2913 (nx15286z55), .px3341 (
                     nx5589z110), .px3342 (nx5589z111), .px3332 (nx5589z106), .px3333 (
                     nx5589z107), .px2894 (nx15286z56), .px2896 (nx15286z57), .px2897 (
                     nx15286z58), .px2898 (nx15286z59), .px2884 (nx15286z60), .px2886 (
                     nx15286z61), .px2887 (nx15286z62), .px2890 (nx15286z63), .px3421 (
                     nx5589z82), .px3422 (nx5589z83), .px3460 (nx5589z11), .px3353 (
                     nx5589z114), .px3354 (nx5589z115), .px3405 (nx5589z53), .px3406 (
                     nx5589z54), .\p_key_samp(4)   (\key_samp(4)  ), .px3392 (
                     nx5589z76), .px3403 (nx5589z77), .px2793 (nx15286z64), .px2794 (
                     nx15286z65), .px2796 (nx15286z66), .px2797 (nx15286z67), .\p_key_samp(45)   (
                     \key_samp(45)  ), .px3307 (nx5589z116), .px3308 (nx5589z117
                     ), .px3335 (nx5589z36), .px2835 (nx15286z68), .px3408 (
                     nx5589z46), .px3338 (nx5589z43), .px2763 (nx15286z69), .px2760 (
                     nx15286z70), .px2892 (nx15286z71), .px2870 (nx15286z72), .px2926 (
                     nx15286z73), .px2773 (nx15286z74), .px2777 (nx15286z75), .px2780 (
                     nx15286z76), .px3304 (nx5589z104), .px3305 (nx5589z105), .px2841 (
                     nx15286z77), .px2866 (nx15286z78), .px2821 (nx15286z79), .px2823 (
                     nx15286z80), .px3359 (nx5589z69), .\p_key_samp(13)   (
                     \key_samp(13)  ), .px3504 (nx5589z94), .px3723 (nx5589z95)
                     , .px3315 (nx5589z100), .px3316 (nx5589z101), .px3321 (
                     nx5589z102), .px3322 (nx5589z103), .px2803 (nx15286z81), .px2810 (
                     nx15286z82), .px2812 (nx15286z83), .\p_key_samp(6)   (
                     \key_samp(6)  ), .px2801 (nx15286z84), .px2867 (nx15286z85)
                     , .px2827 (nx15286z86), .px2698 (nx15286z87), .px2702 (
                     nx15286z88), .px2703 (nx15286z89), .\p_key_samp(61)   (
                     \key_samp(61)  ), .px2733 (nx15286z90), .px2741 (nx15286z91
                     ), .px2723 (nx15286z92), .px2729 (nx15286z93), .px2711 (
                     nx15286z94), .px2712 (nx15286z95), .px2764 (nx15286z96), .px2751 (
                     nx15286z97), .\p_key_samp(10)   (\key_samp(10)  ), .\p_key_samp(46)   (
                     \key_samp(46)  ), .px2680 (nx15286z98), .px2682 (nx15286z99
                     ), .px2683 (nx15286z100), .px2694 (nx15286z101), .\p_key_samp(21)   (
                     \key_samp(21)  ), .\p_key_samp(12)   (\key_samp(12)  ), .\p_key_samp(5)   (
                     \key_samp(5)  ), .\p_key_samp(7)   (\key_samp(7)  ), .px2765 (
                     nx15286z102), .px2719 (nx15286z103), .px2709 (nx15286z104)
                     , .px2731 (nx15286z105), .\p_key_samp(49)   (\key_samp(49)  
                     ), .px2642 (nx15286z106), .px2643 (nx15286z107), .px2644 (
                     nx15286z108), .px2646 (nx15286z109), .px2618 (nx15286z110)
                     , .px2621 (nx15286z111), .px2622 (nx15286z112), .px2623 (
                     nx15286z113), .\p_key_samp(39)   (\key_samp(39)  ), .\p_key_samp(47)   (
                     \key_samp(47)  ), .\p_key_samp(28)   (\key_samp(28)  ), .px2654 (
                     nx15286z114), .px2656 (nx15286z115), .px2658 (nx15286z116)
                     , .px2664 (nx15286z117), .\p_key_samp(23)   (\key_samp(23)  
                     ), .px2630 (nx15286z118), .px2634 (nx15286z119), .px2637 (
                     nx15286z120), .px2638 (nx15286z121), .\p_key_samp(22)   (
                     \key_samp(22)  ), .\p_key_samp(54)   (\key_samp(54)  ), .\p_key_samp(37)   (
                     \key_samp(37)  ), .px2668 (nx15286z122), .px2670 (
                     nx15286z123), .px2669 (nx15286z124), .px2672 (nx15286z125)
                     , .px2605 (nx15286z126), .px2606 (nx15286z127), .px2607 (
                     nx15286z128), .px2608 (nx15286z129), .px3007 (nx5589z273), 
                     .\p_key_samp(14)   (\key_samp(14)  ), .\p_key_samp(63)   (
                     \key_samp(63)  ), .\p_key_samp(30)   (\key_samp(30)  ), .\p_key_samp(53)   (
                     \key_samp(53)  ), .\p_key_samp(31)   (\key_samp(31)  ), .px2514 (
                     nx15286z130), .px2507 (nx15286z131), .\p_key_samp(29)   (
                     \key_samp(29)  ), .\p_key_samp(20)   (\key_samp(20)  ), .px3036 (
                     nx5589z278), .\p_key_samp(62)   (\key_samp(62)  ), .\p_key_samp(38)   (
                     \key_samp(38)  ), .\p_key_samp(55)   (\key_samp(55)  ), .px2497 (
                     nx15286z132), .\p_key_samp(19)   (\key_samp(19)  ), .\p_key_samp(52)   (
                     \key_samp(52)  ), .px3052 (nx5589z283), .\p_key_samp(59)   (
                     \key_samp(59)  ), .\p_key_samp(34)   (\key_samp(34)  ), .\p_key_samp(2)   (
                     \key_samp(2)  ), .\p_key_samp(17)   (\key_samp(17)  ), .\p_key_samp(26)   (
                     \key_samp(26)  ), .px2585 (nx15286z133), .px2591 (
                     nx15286z134), .px2587 (nx15286z135), .px2593 (nx15286z136)
                     , .\p_key_samp(51)   (\key_samp(51)  ), .\p_key_samp(3)   (
                     \key_samp(3)  ), .\p_key_samp(33)   (\key_samp(33)  ), .\p_key_samp(9)   (
                     \key_samp(9)  ), .px2628 (nx15286z137), .px2640 (
                     nx15286z138), .px2678 (nx15286z139), .px2706 (nx15286z140)
                     , .\p_key_samp(27)   (\key_samp(27)  ), .\p_key_samp(35)   (
                     \key_samp(35)  ), .\p_key_samp(58)   (\key_samp(58)  ), .px2570 (
                     nx15286z141), .px2569 (nx15286z142), .px2566 (nx15286z143)
                     , .px2563 (nx15286z144), .\p_key_samp(36)   (\key_samp(36)  
                     ), .px2573 (nx15286z145), .px2575 (nx15286z146), .px2579 (
                     nx15286z147), .px2582 (nx15286z148), .\p_key_samp(18)   (
                     \key_samp(18)  ), .px2601 (nx15286z149), .px2611 (
                     nx15286z150), .px2613 (nx15286z151), .px2615 (nx15286z152)
                     , .\p_key_samp(41)   (\key_samp(41)  ), .px2551 (
                     nx15286z153), .px2555 (nx15286z154), .px2557 (nx15286z155)
                     , .px2558 (nx15286z156), .\p_key_samp(60)   (\key_samp(60)  
                     ), .\p_key_samp(25)   (\key_samp(25)  ), .\p_key_samp(42)   (
                     \key_samp(42)  ), .\p_key_samp(1)   (\key_samp(1)  ), .\p_key_samp(11)   (
                     \key_samp(11)  ), .px2528 (nx15286z157), .px2523 (
                     nx15286z158), .px2522 (nx15286z159), .px2521 (nx15286z160)
                     , .\p_key_samp(57)   (\key_samp(57)  ), .px2537 (
                     nx15286z161), .px2534 (nx15286z162), .px2533 (nx15286z163)
                     , .px2538 (nx15286z164), .\p_key_samp(43)   (\key_samp(43)  
                     ), .px2708 (nx5589z244), .px2869 (nx5589z245), .px3058 (
                     nx5589z246), .px3281 (nx5589z247), .px3503 (nx5589z248), .px2432 (
                     nx18561z1), .px2707 (nx5589z194), .px2868 (nx5589z195), .px3057 (
                     nx5589z196), .px3221 (nx5589z197), .px3222 (nx5589z198), .px2431 (
                     nx20555z1), .px2430 (nx59360z1), .px2429 (nx56367z1), .px2576 (
                     nx5589z239), .px2742 (nx5589z240), .px2891 (nx5589z241), .px3092 (
                     nx5589z242), .px3093 (nx5589z243), .px2428 (nx43404z1), .px2588 (
                     nx5589z219), .px2768 (nx5589z220), .px2941 (nx5589z221), .px3151 (
                     nx5589z222), .px3152 (nx5589z223), .px2427 (nx30441z1), .px2426 (
                     nx19472z1), .px2425 (nx15484z1), .px2592 (nx5589z199), .px2786 (
                     nx5589z200), .px2945 (nx5589z201), .px3160 (nx5589z202), .px3161 (
                     nx5589z203), .px2424 (nx1800z1), .px2641 (nx5589z189), .px2828 (
                     nx5589z190), .px2953 (nx5589z191), .px3187 (nx5589z192), .px3202 (
                     nx5589z193), .px2423 (nx4793z1), .px2422 (nx48391z1), .px2421 (
                     nx54373z1), .px2420 (nx14573z1), .px2629 (nx5589z209), .px2802 (
                     nx5589z210), .px3017 (nx5589z211), .px3170 (nx5589z212), .px3185 (
                     nx5589z213), .px2419 (nx32435z1), .px2418 (nx17478z1), .px2556 (
                     nx5589z259), .px2730 (nx5589z260), .px2899 (nx5589z261), .px3068 (
                     nx5589z262), .px3069 (nx5589z263), .px2417 (nx16567z1), .px2602 (
                     nx5589z229), .px2748 (nx5589z230), .px2914 (nx5589z231), .px3119 (
                     nx5589z232), .px3120 (nx5589z233), .px2416 (nx6787z1), .px2415 (
                     nx52379z1), .px2594 (nx5589z214), .px2772 (nx5589z215), .px2929 (
                     nx5589z216), .px3138 (nx5589z217), .px3149 (nx5589z218), .px2414 (
                     nx22549z1), .px2413 (nx28447z1), .px2614 (nx5589z264), .px2752 (
                     nx5589z265), .px2909 (nx5589z266), .px3112 (nx5589z267), .px3113 (
                     nx5589z268), .px2412 (nx37422z1), .px2586 (nx5589z224), .px2770 (
                     nx5589z225), .px2943 (nx5589z226), .px3154 (nx5589z227), .px3155 (
                     nx5589z228), .px2411 (nx39416z1), .px2410 (nx26453z1), .px2409 (
                     nx23460z1), .px2552 (nx5589z249), .px2728 (nx5589z250), .px2895 (
                     nx5589z251), .px3073 (nx5589z252), .px3074 (nx5589z253), .px2408 (
                     nx65342z1), .px2574 (nx5589z234), .px2734 (nx5589z235), .px2885 (
                     nx5589z236), .px3095 (nx5589z237), .px3096 (nx5589z238), .px2407 (
                     nx34429z1), .px2406 (nx50385z1), .px2405 (nx63348z1), .px2612 (
                     nx5589z254), .px2746 (nx5589z255), .px2907 (nx5589z256), .px3109 (
                     nx5589z257), .px3110 (nx5589z258), .px2404 (nx45398z1), .px2403 (
                     nx21466z1), .px2402 (nx61354z1), .px2679 (nx5589z204), .px2790 (
                     nx5589z205), .px2985 (nx5589z206), .px3245 (nx5589z207), .px3280 (
                     nx5589z208), .px2401 (nx41410z1), .px2671 (nx5589z138), .px2855 (
                     nx5589z139), .px3010 (nx5589z140), .px3216 (nx5589z141), .px3217 (
                     nx5589z142), .px2400 (nx63706z1), .px2639 (nx5589z182), .px2807 (
                     nx5589z183), .px3022 (nx5589z184), .px3172 (nx5589z185), .px3173 (
                     nx5589z186), .px2399 (nx164z1), .px2665 (nx5589z167), .px2820 (
                     nx5589z168), .px2973 (nx5589z169), .px3232 (nx5589z170), .px3233 (
                     nx5589z171), .px2398 (nx3157z1), .px2766 (nx5589z123), .px2927 (
                     nx5589z124), .px3136 (nx5589z125), .px3330 (nx5589z126), .px3349 (
                     nx5589z127), .px2397 (nx5151z1), .px2396 (nx7145z1), .px2395 (
                     nx9139z1), .px2394 (nx11133z1), .px2393 (nx14126z1), .px2392 (
                     nx16120z1), .px2391 (nx18114z1), .px2390 (nx20108z1), .px2389 (
                     nx22102z1), .px2720 (nx5589z133), .px2893 (nx5589z134), .px3060 (
                     nx5589z135), .px3296 (nx5589z136), .px3311 (nx5589z137), .px2388 (
                     nx25095z1), .px2647 (nx5589z145), .px2832 (nx5589z146), .px3054 (
                     nx5589z147), .px3197 (nx5589z148), .px3198 (nx5589z149), .px2387 (
                     nx27089z1), .px2655 (nx5589z177), .px2818 (nx5589z178), .px2970 (
                     nx5589z179), .px3229 (nx5589z180), .px3230 (nx5589z181), .px2386 (
                     nx29083z1), .px2695 (nx5589z157), .px2798 (nx5589z158), .px2997 (
                     nx5589z159), .px3278 (nx5589z160), .px3279 (nx5589z161), .px2385 (
                     nx31077z1), .px2710 (nx5589z128), .px2871 (nx5589z129), .px3077 (
                     nx5589z130), .px3283 (nx5589z131), .px3294 (nx5589z132), .px2384 (
                     nx33071z1), .px2508 (nx5589z274), .px2645 (nx5589z275), .px2836 (
                     nx5589z276), .px3035 (nx5589z277), .px3191 (nx5589z150), .px3192 (
                     nx5589z151), .px2383 (nx36064z1), .px2657 (nx5589z172), .px2822 (
                     nx5589z173), .px2967 (nx5589z174), .px3226 (nx5589z175), .px3227 (
                     nx5589z176), .px2382 (nx38058z1), .px2681 (nx5589z162), .px2795 (
                     nx5589z163), .px2987 (nx5589z164), .px3261 (nx5589z165), .px3262 (
                     nx5589z166), .px2381 (nx40052z1), .px2380 (nx42046z1), .px2379 (
                     nx44040z1), .px2378 (nx47033z1), .px2377 (nx49027z1), .px2376 (
                     nx51021z1), .px2375 (nx53015z1), .px2374 (nx55009z1), .px2373 (
                     nx65314z1), .px2732 (nx5589z118), .px2881 (nx5589z119), .px3090 (
                     nx5589z120), .px3313 (nx5589z121), .px3328 (nx5589z122), .px2372 (
                     nx1772z1), .px2520 (nx5589z269), .px2673 (nx5589z270), .px2857 (
                     nx5589z271), .px3006 (nx5589z272), .px3206 (nx5589z143), .px3207 (
                     nx5589z144), .px2371 (nx3766z1), .px2498 (nx5589z279), .px2631 (
                     nx5589z280), .px2811 (nx5589z281), .px3041 (nx5589z282), .px3183 (
                     nx5589z187), .px3184 (nx5589z188), .px2370 (nx5760z1), .px2659 (
                     nx5589z152), .px2824 (nx5589z153), .px2982 (nx5589z154), .px3235 (
                     nx5589z155), .px3236 (nx5589z156), .px2369 (nx7754z1), .p_nbus_data_in_int (
                     {data_in_int[0],data_in_int[1],data_in_int[2],
                     data_in_int[3],data_in_int[4],data_in_int[5],data_in_int[6]
                     ,data_in_int[7],data_in_int[8],data_in_int[9],
                     data_in_int[10],data_in_int[11],data_in_int[12],
                     data_in_int[13],data_in_int[14],data_in_int[15],
                     data_in_int[16],data_in_int[17],data_in_int[18],
                     data_in_int[19],data_in_int[20],data_in_int[21],
                     data_in_int[22],data_in_int[23],data_in_int[24],
                     data_in_int[25],data_in_int[26],data_in_int[27],
                     data_in_int[28],data_in_int[29],data_in_int[30],
                     data_in_int[31],data_in_int[32],data_in_int[33],
                     data_in_int[34],data_in_int[35],data_in_int[36],
                     data_in_int[37],data_in_int[38],data_in_int[39],
                     data_in_int[40],data_in_int[41],data_in_int[42],
                     data_in_int[43],data_in_int[44],data_in_int[45],
                     data_in_int[46],data_in_int[47],data_in_int[48],
                     data_in_int[49],data_in_int[50],data_in_int[51],
                     data_in_int[52],data_in_int[53],data_in_int[54],
                     data_in_int[55],data_in_int[56],data_in_int[57],
                     data_in_int[58],data_in_int[59],data_in_int[60],
                     data_in_int[61],data_in_int[62],data_in_int[63]}), .p_nbus_plaintext (
                     {\plaintext(5)  }), .\p_plaintext(37)   (\plaintext(37)  )
                     , .\p_plaintext(39)   (\plaintext(39)  ), .p_reset_int (
                     reset_int), .p_load_int (load_int), .p_clk_int (clk_int), .\p_plaintext(63)   (
                     \plaintext(63)  )) ;
    input_register_1 i_key_samp (.\p_plaintext(5)   (\plaintext(5)  ), .px3923 (
                     nx15286z3), .px3872 (nx15286z2), .\p_plaintext(63)   (
                     \plaintext(63)  ), .px3870 (nx15286z1), .px3745 (nx5589z1)
                     , .\p_plaintext(37)   (\plaintext(37)  ), .px3744 (
                     nx15286z5), .px3781 (nx5589z2), .\p_plaintext(39)   (
                     \plaintext(39)  ), .px3697 (nx15286z4), .px3089 (nx15286z11
                     ), .px3076 (nx15286z13), .px3059 (nx15286z12), .px3056 (
                     nx15286z39), .px3635 (nx5589z3), .px3636 (nx5589z4), .px3053 (
                     nx15286z31), .px3040 (nx15286z30), .px3034 (nx15286z29), .px3021 (
                     nx15286z28), .px3016 (nx15286z38), .px3752 (nx5589z5), .px3761 (
                     nx5589z6), .px3015 (nx15286z23), .px3726 (nx5589z7), .px3737 (
                     nx5589z8), .px3008 (nx15286z22), .px3005 (nx15286z21), .px3739 (
                     nx5589z9), .px3750 (nx5589z10), .px2999 (nx15286z10), .px2996 (
                     nx15286z9), .px2986 (nx15286z8), .px2984 (nx15286z37), .px2981 (
                     nx15286z27), .px3460 (nx5589z11), .px3705 (nx5589z12), .px3714 (
                     nx5589z13), .px2972 (nx15286z26), .px2969 (nx15286z25), .px2966 (
                     nx15286z24), .px3638 (nx5589z14), .px3639 (nx5589z15), .px2963 (
                     nx15286z7), .px3483 (nx5589z16), .px3674 (nx5589z17), .px3675 (
                     nx5589z18), .px2959 (nx15286z6), .px2952 (nx15286z36), .px2944 (
                     nx15286z33), .px2942 (nx15286z34), .px2940 (nx15286z35), .px3448 (
                     nx5589z19), .px3688 (nx5589z20), .px3689 (nx5589z21), .px2939 (
                     nx15286z20), .px3716 (nx5589z22), .px3717 (nx5589z23), .px2935 (
                     nx15286z19), .px3626 (nx5589z24), .px3627 (nx5589z25), .px2934 (
                     nx15286z18), .px3623 (nx5589z26), .px3624 (nx5589z27), .px2933 (
                     nx15286z17), .px2928 (nx15286z32), .px2926 (nx15286z73), .px3702 (
                     nx5589z28), .px3703 (nx5589z29), .px2925 (nx15286z15), .px3657 (
                     nx5589z30), .px3658 (nx5589z31), .px2924 (nx15286z16), .px3665 (
                     nx5589z32), .px3666 (nx5589z33), .px2921 (nx15286z14), .px2913 (
                     nx15286z55), .px2912 (nx15286z52), .px2908 (nx15286z53), .px2906 (
                     nx15286z54), .px2898 (nx15286z59), .px3584 (nx5589z34), .px3585 (
                     nx5589z35), .px2897 (nx15286z58), .px3335 (nx5589z36), .px3590 (
                     nx5589z37), .px3591 (nx5589z38), .px2896 (nx15286z57), .px2894 (
                     nx15286z56), .px2892 (nx15286z71), .px2890 (nx15286z63), .px3649 (
                     nx5589z39), .px3650 (nx5589z40), .px2887 (nx15286z62), .px3632 (
                     nx5589z41), .px3647 (nx5589z42), .px2886 (nx15286z61), .px2884 (
                     nx15286z60), .px3338 (nx5589z43), .px3546 (nx5589z44), .px3547 (
                     nx5589z45), .px2879 (nx15286z51), .px3408 (nx5589z46), .px3652 (
                     nx5589z47), .px3667 (nx5589z48), .px2878 (nx15286z50), .px3615 (
                     nx5589z49), .px3630 (nx5589z50), .px2877 (nx15286z49), .px3543 (
                     nx5589z51), .px3544 (nx5589z52), .px2872 (nx15286z48), .px2870 (
                     nx15286z72), .px3405 (nx5589z53), .px3406 (nx5589z54), .px2867 (
                     nx15286z85), .px3523 (nx5589z55), .px3534 (nx5589z56), .px2866 (
                     nx15286z78), .px3596 (nx5589z57), .px3607 (nx5589z58), .px2865 (
                     nx15286z40), .px3587 (nx5589z59), .px3588 (nx5589z60), .px2860 (
                     nx15286z43), .px3559 (nx5589z61), .px3560 (nx5589z62), .px2859 (
                     nx15286z41), .px3562 (nx5589z63), .px3563 (nx5589z64), .px2858 (
                     nx15286z42), .px3514 (nx5589z65), .px3515 (nx5589z66), .px2847 (
                     nx15286z47), .px3511 (nx5589z67), .px3512 (nx5589z68), .px2846 (
                     nx15286z46), .px3359 (nx5589z69), .px3565 (nx5589z70), .px3576 (
                     nx5589z71), .px2845 (nx15286z45), .px3724 (nx5589z72), .px3886 (
                     nx5589z73), .px2844 (nx15286z44), .px3582 (nx5589z74), .px3611 (
                     nx5589z75), .px2841 (nx15286z77), .px2835 (nx15286z68), .px3392 (
                     nx5589z76), .px3403 (nx5589z77), .px2827 (nx15286z86), .px2823 (
                     nx15286z80), .px2821 (nx15286z79), .px3436 (nx5589z78), .px3437 (
                     nx5589z79), .px2812 (nx15286z83), .px2810 (nx15286z82), .px3442 (
                     nx5589z80), .px3443 (nx5589z81), .px2803 (nx15286z81), .px2801 (
                     nx15286z84), .px3421 (nx5589z82), .px3422 (nx5589z83), .px2797 (
                     nx15286z67), .px3506 (nx5589z84), .px3521 (nx5589z85), .px2796 (
                     nx15286z66), .px2794 (nx15286z65), .px3536 (nx5589z86), .px3551 (
                     nx5589z87), .px2793 (nx15286z64), .px3439 (nx5589z88), .px3440 (
                     nx5589z89), .px2780 (nx15286z76), .px3454 (nx5589z90), .px3455 (
                     nx5589z91), .px2777 (nx15286z75), .px3433 (nx5589z92), .px3434 (
                     nx5589z93), .px2773 (nx15286z74), .px2765 (nx15286z102), .px3504 (
                     nx5589z94), .px3723 (nx5589z95), .px2764 (nx15286z96), .px3451 (
                     nx5589z96), .px3452 (nx5589z97), .px2763 (nx15286z69), .px3410 (
                     nx5589z98), .px3411 (nx5589z99), .px2760 (nx15286z70), .px2751 (
                     nx15286z97), .px3315 (nx5589z100), .px3316 (nx5589z101), .px2741 (
                     nx15286z91), .px3321 (nx5589z102), .px3322 (nx5589z103), .px2733 (
                     nx15286z90), .px2731 (nx15286z105), .px3304 (nx5589z104), .px3305 (
                     nx5589z105), .px2729 (nx15286z93), .px3332 (nx5589z106), .px3333 (
                     nx5589z107), .px2723 (nx15286z92), .px2719 (nx15286z103), .px3425 (
                     nx5589z108), .px3444 (nx5589z109), .px2712 (nx15286z95), .px3341 (
                     nx5589z110), .px3342 (nx5589z111), .px2711 (nx15286z94), .px2709 (
                     nx15286z104), .px2706 (nx15286z140), .px3373 (nx5589z112), 
                     .px3374 (nx5589z113), .px2703 (nx15286z89), .px3353 (
                     nx5589z114), .px3354 (nx5589z115), .px2702 (nx15286z88), .px3307 (
                     nx5589z116), .px3308 (nx5589z117), .px2698 (nx15286z87), .px2694 (
                     nx15286z101), .px2732 (nx5589z118), .px2881 (nx5589z119), .px3090 (
                     nx5589z120), .px3313 (nx5589z121), .px3328 (nx5589z122), .px2683 (
                     nx15286z100), .px2766 (nx5589z123), .px2927 (nx5589z124), .px3136 (
                     nx5589z125), .px3330 (nx5589z126), .px3349 (nx5589z127), .px2682 (
                     nx15286z99), .px2680 (nx15286z98), .px2678 (nx15286z139), .px2672 (
                     nx15286z125), .px2670 (nx15286z123), .px2710 (nx5589z128), 
                     .px2871 (nx5589z129), .px3077 (nx5589z130), .px3283 (
                     nx5589z131), .px3294 (nx5589z132), .px2669 (nx15286z124), .px2720 (
                     nx5589z133), .px2893 (nx5589z134), .px3060 (nx5589z135), .px3296 (
                     nx5589z136), .px3311 (nx5589z137), .px2668 (nx15286z122), .px2664 (
                     nx15286z117), .px2658 (nx15286z116), .px2656 (nx15286z115)
                     , .px2654 (nx15286z114), .px2646 (nx15286z109), .px2644 (
                     nx15286z108), .px2671 (nx5589z138), .px2855 (nx5589z139), .px3010 (
                     nx5589z140), .px3216 (nx5589z141), .px3217 (nx5589z142), .px2643 (
                     nx15286z107), .px3206 (nx5589z143), .px3207 (nx5589z144), .px2642 (
                     nx15286z106), .px2640 (nx15286z138), .px2638 (nx15286z121)
                     , .px2647 (nx5589z145), .px2832 (nx5589z146), .px3054 (
                     nx5589z147), .px3197 (nx5589z148), .px3198 (nx5589z149), .px2637 (
                     nx15286z120), .px3191 (nx5589z150), .px3192 (nx5589z151), .px2634 (
                     nx15286z119), .px2630 (nx15286z118), .px2628 (nx15286z137)
                     , .px2659 (nx5589z152), .px2824 (nx5589z153), .px2982 (
                     nx5589z154), .px3235 (nx5589z155), .px3236 (nx5589z156), .px2623 (
                     nx15286z113), .px2695 (nx5589z157), .px2798 (nx5589z158), .px2997 (
                     nx5589z159), .px3278 (nx5589z160), .px3279 (nx5589z161), .px2622 (
                     nx15286z112), .px2681 (nx5589z162), .px2795 (nx5589z163), .px2987 (
                     nx5589z164), .px3261 (nx5589z165), .px3262 (nx5589z166), .px2621 (
                     nx15286z111), .px2665 (nx5589z167), .px2820 (nx5589z168), .px2973 (
                     nx5589z169), .px3232 (nx5589z170), .px3233 (nx5589z171), .px2618 (
                     nx15286z110), .px2615 (nx15286z152), .px2613 (nx15286z151)
                     , .px2611 (nx15286z150), .px2657 (nx5589z172), .px2822 (
                     nx5589z173), .px2967 (nx5589z174), .px3226 (nx5589z175), .px3227 (
                     nx5589z176), .px2608 (nx15286z129), .px2655 (nx5589z177), .px2818 (
                     nx5589z178), .px2970 (nx5589z179), .px3229 (nx5589z180), .px3230 (
                     nx5589z181), .px2607 (nx15286z128), .px2639 (nx5589z182), .px2807 (
                     nx5589z183), .px3022 (nx5589z184), .px3172 (nx5589z185), .px3173 (
                     nx5589z186), .px2606 (nx15286z127), .px3183 (nx5589z187), .px3184 (
                     nx5589z188), .px2605 (nx15286z126), .px2601 (nx15286z149), 
                     .px2593 (nx15286z136), .px2591 (nx15286z134), .px2587 (
                     nx15286z135), .px2585 (nx15286z133), .px2641 (nx5589z189), 
                     .px2828 (nx5589z190), .px2953 (nx5589z191), .px3187 (
                     nx5589z192), .px3202 (nx5589z193), .px2582 (nx15286z148), .px2707 (
                     nx5589z194), .px2868 (nx5589z195), .px3057 (nx5589z196), .px3221 (
                     nx5589z197), .px3222 (nx5589z198), .px2579 (nx15286z147), .px2575 (
                     nx15286z146), .px2573 (nx15286z145), .px2592 (nx5589z199), 
                     .px2786 (nx5589z200), .px2945 (nx5589z201), .px3160 (
                     nx5589z202), .px3161 (nx5589z203), .px2570 (nx15286z141), .px2679 (
                     nx5589z204), .px2790 (nx5589z205), .px2985 (nx5589z206), .px3245 (
                     nx5589z207), .px3280 (nx5589z208), .px2569 (nx15286z142), .px2629 (
                     nx5589z209), .px2802 (nx5589z210), .px3017 (nx5589z211), .px3170 (
                     nx5589z212), .px3185 (nx5589z213), .px2566 (nx15286z143), .px2594 (
                     nx5589z214), .px2772 (nx5589z215), .px2929 (nx5589z216), .px3138 (
                     nx5589z217), .px3149 (nx5589z218), .px2563 (nx15286z144), .px2588 (
                     nx5589z219), .px2768 (nx5589z220), .px2941 (nx5589z221), .px3151 (
                     nx5589z222), .px3152 (nx5589z223), .px2558 (nx15286z156), .px2586 (
                     nx5589z224), .px2770 (nx5589z225), .px2943 (nx5589z226), .px3154 (
                     nx5589z227), .px3155 (nx5589z228), .px2557 (nx15286z155), .px2555 (
                     nx15286z154), .px2551 (nx15286z153), .px2602 (nx5589z229), 
                     .px2748 (nx5589z230), .px2914 (nx5589z231), .px3119 (
                     nx5589z232), .px3120 (nx5589z233), .px2538 (nx15286z164), .px2574 (
                     nx5589z234), .px2734 (nx5589z235), .px2885 (nx5589z236), .px3095 (
                     nx5589z237), .px3096 (nx5589z238), .px2537 (nx15286z161), .px2576 (
                     nx5589z239), .px2742 (nx5589z240), .px2891 (nx5589z241), .px3092 (
                     nx5589z242), .px3093 (nx5589z243), .px2534 (nx15286z162), .px2708 (
                     nx5589z244), .px2869 (nx5589z245), .px3058 (nx5589z246), .px3281 (
                     nx5589z247), .px3503 (nx5589z248), .px2533 (nx15286z163), .px2552 (
                     nx5589z249), .px2728 (nx5589z250), .px2895 (nx5589z251), .px3073 (
                     nx5589z252), .px3074 (nx5589z253), .px2528 (nx15286z157), .px2612 (
                     nx5589z254), .px2746 (nx5589z255), .px2907 (nx5589z256), .px3109 (
                     nx5589z257), .px3110 (nx5589z258), .px2523 (nx15286z158), .px2556 (
                     nx5589z259), .px2730 (nx5589z260), .px2899 (nx5589z261), .px3068 (
                     nx5589z262), .px3069 (nx5589z263), .px2522 (nx15286z159), .px2614 (
                     nx5589z264), .px2752 (nx5589z265), .px2909 (nx5589z266), .px3112 (
                     nx5589z267), .px3113 (nx5589z268), .px2521 (nx15286z160), .px2520 (
                     nx5589z269), .px2673 (nx5589z270), .px2857 (nx5589z271), .px3006 (
                     nx5589z272), .px3007 (nx5589z273), .px2514 (nx15286z130), .px2508 (
                     nx5589z274), .px2645 (nx5589z275), .px2836 (nx5589z276), .px3035 (
                     nx5589z277), .px3036 (nx5589z278), .px2507 (nx15286z131), .px2498 (
                     nx5589z279), .px2631 (nx5589z280), .px2811 (nx5589z281), .px3041 (
                     nx5589z282), .px3052 (nx5589z283), .px2497 (nx15286z132), .p_nbus_key_in_int (
                     {key_in_int[8],key_in_int[9],key_in_int[10],key_in_int[11],
                     key_in_int[12],key_in_int[13],key_in_int[14],key_in_int[15]
                     ,key_in_int[16],key_in_int[17],key_in_int[18],
                     key_in_int[19],key_in_int[20],key_in_int[21],key_in_int[22]
                     ,key_in_int[23],key_in_int[24],key_in_int[25],
                     key_in_int[26],key_in_int[27],key_in_int[28],key_in_int[29]
                     ,key_in_int[30],key_in_int[31],key_in_int[32],
                     key_in_int[33],key_in_int[34],key_in_int[35],key_in_int[36]
                     ,key_in_int[37],key_in_int[38],key_in_int[39],
                     key_in_int[40],key_in_int[41],key_in_int[42],key_in_int[43]
                     ,key_in_int[44],key_in_int[45],key_in_int[46],
                     key_in_int[47],key_in_int[48],key_in_int[49],key_in_int[50]
                     ,key_in_int[51],key_in_int[52],key_in_int[53],
                     key_in_int[54],key_in_int[55],key_in_int[56],key_in_int[57]
                     ,key_in_int[58],key_in_int[59],key_in_int[60],
                     key_in_int[61],key_in_int[62],key_in_int[63]}), .\p_key_samp(1)   (
                     \key_samp(1)  ), .\p_key_samp(2)   (\key_samp(2)  ), .\p_key_samp(3)   (
                     \key_samp(3)  ), .\p_key_samp(4)   (\key_samp(4)  ), .\p_key_samp(5)   (
                     \key_samp(5)  ), .\p_key_samp(6)   (\key_samp(6)  ), .\p_key_samp(7)   (
                     \key_samp(7)  ), .\p_key_samp(9)   (\key_samp(9)  ), .\p_key_samp(10)   (
                     \key_samp(10)  ), .\p_key_samp(11)   (\key_samp(11)  ), .\p_key_samp(12)   (
                     \key_samp(12)  ), .\p_key_samp(13)   (\key_samp(13)  ), .\p_key_samp(14)   (
                     \key_samp(14)  ), .\p_key_samp(15)   (\key_samp(15)  ), .\p_key_samp(17)   (
                     \key_samp(17)  ), .\p_key_samp(18)   (\key_samp(18)  ), .\p_key_samp(19)   (
                     \key_samp(19)  ), .\p_key_samp(20)   (\key_samp(20)  ), .\p_key_samp(21)   (
                     \key_samp(21)  ), .\p_key_samp(22)   (\key_samp(22)  ), .\p_key_samp(23)   (
                     \key_samp(23)  ), .\p_key_samp(25)   (\key_samp(25)  ), .\p_key_samp(26)   (
                     \key_samp(26)  ), .\p_key_samp(27)   (\key_samp(27)  ), .\p_key_samp(28)   (
                     \key_samp(28)  ), .\p_key_samp(29)   (\key_samp(29)  ), .\p_key_samp(30)   (
                     \key_samp(30)  ), .\p_key_samp(31)   (\key_samp(31)  ), .\p_key_samp(33)   (
                     \key_samp(33)  ), .\p_key_samp(34)   (\key_samp(34)  ), .\p_key_samp(35)   (
                     \key_samp(35)  ), .\p_key_samp(36)   (\key_samp(36)  ), .\p_key_samp(37)   (
                     \key_samp(37)  ), .\p_key_samp(38)   (\key_samp(38)  ), .\p_key_samp(39)   (
                     \key_samp(39)  ), .\p_key_samp(41)   (\key_samp(41)  ), .\p_key_samp(42)   (
                     \key_samp(42)  ), .\p_key_samp(43)   (\key_samp(43)  ), .\p_key_samp(44)   (
                     \key_samp(44)  ), .\p_key_samp(45)   (\key_samp(45)  ), .\p_key_samp(46)   (
                     \key_samp(46)  ), .\p_key_samp(47)   (\key_samp(47)  ), .\p_key_samp(49)   (
                     \key_samp(49)  ), .\p_key_samp(50)   (\key_samp(50)  ), .\p_key_samp(51)   (
                     \key_samp(51)  ), .\p_key_samp(52)   (\key_samp(52)  ), .\p_key_samp(53)   (
                     \key_samp(53)  ), .\p_key_samp(54)   (\key_samp(54)  ), .\p_key_samp(55)   (
                     \key_samp(55)  ), .\p_key_samp(57)   (\key_samp(57)  ), .\p_key_samp(58)   (
                     \key_samp(58)  ), .\p_key_samp(59)   (\key_samp(59)  ), .\p_key_samp(60)   (
                     \key_samp(60)  ), .\p_key_samp(61)   (\key_samp(61)  ), .\p_key_samp(62)   (
                     \key_samp(62)  ), .p_reset_int (reset_int), .p_load_int (
                     load_int), .p_clk_int (clk_int), .\p_key_samp(63)   (
                     \key_samp(63)  )) ;
    BUFGP clk_ibuf (.O (clk_int), .I (clk)) ;
    VCC \reg_data_out(4)_I22_FD_PWR  (.P (nx4)) ;
    FDRE \reg_data_out(4)  (.Q (data_out_1_0[4]), .C (clk_int), .CE (nx4), .D (
         nx18561z1), .R (reset_int)) ;
    FDRE \reg_data_out(2)  (.Q (data_out_1_0[2]), .C (clk_int), .CE (nx4), .D (
         nx20555z1), .R (reset_int)) ;
    FDRE \reg_data_out(50)  (.Q (data_out_1_0[50]), .C (clk_int), .CE (nx4), .D (
         nx59360z1), .R (reset_int)) ;
    FDRE \reg_data_out(48)  (.Q (data_out_1_0[48]), .C (clk_int), .CE (nx4), .D (
         nx56367z1), .R (reset_int)) ;
    FDRE \reg_data_out(36)  (.Q (data_out_1_0[36]), .C (clk_int), .CE (nx4), .D (
         nx43404z1), .R (reset_int)) ;
    FDRE \reg_data_out(24)  (.Q (data_out_1_0[24]), .C (clk_int), .CE (nx4), .D (
         nx30441z1), .R (reset_int)) ;
    FDRE \reg_data_out(14)  (.Q (data_out_1_0[14]), .C (clk_int), .CE (nx4), .D (
         nx19472z1), .R (reset_int)) ;
    FDRE \reg_data_out(10)  (.Q (data_out_1_0[10]), .C (clk_int), .CE (nx4), .D (
         nx15484z1), .R (reset_int)) ;
    FDRE \reg_data_out(58)  (.Q (data_out_1_0[58]), .C (clk_int), .CE (nx4), .D (
         nx1800z1), .R (reset_int)) ;
    FDRE \reg_data_out(60)  (.Q (data_out_1_0[60]), .C (clk_int), .CE (nx4), .D (
         nx4793z1), .R (reset_int)) ;
    FDRE \reg_data_out(40)  (.Q (data_out_1_0[40]), .C (clk_int), .CE (nx4), .D (
         nx48391z1), .R (reset_int)) ;
    FDRE \reg_data_out(46)  (.Q (data_out_1_0[46]), .C (clk_int), .CE (nx4), .D (
         nx54373z1), .R (reset_int)) ;
    FDRE \reg_data_out(8)  (.Q (data_out_1_0[8]), .C (clk_int), .CE (nx4), .D (
         nx14573z1), .R (reset_int)) ;
    FDRE \reg_data_out(26)  (.Q (data_out_1_0[26]), .C (clk_int), .CE (nx4), .D (
         nx32435z1), .R (reset_int)) ;
    FDRE \reg_data_out(12)  (.Q (data_out_1_0[12]), .C (clk_int), .CE (nx4), .D (
         nx17478z1), .R (reset_int)) ;
    FDRE \reg_data_out(6)  (.Q (data_out_1_0[6]), .C (clk_int), .CE (nx4), .D (
         nx16567z1), .R (reset_int)) ;
    FDRE \reg_data_out(62)  (.Q (data_out_1_0[62]), .C (clk_int), .CE (nx4), .D (
         nx6787z1), .R (reset_int)) ;
    FDRE \reg_data_out(44)  (.Q (data_out_1_0[44]), .C (clk_int), .CE (nx4), .D (
         nx52379z1), .R (reset_int)) ;
    FDRE \reg_data_out(0)  (.Q (data_out_1_0[0]), .C (clk_int), .CE (nx4), .D (
         nx22549z1), .R (reset_int)) ;
    FDRE \reg_data_out(22)  (.Q (data_out_1_0[22]), .C (clk_int), .CE (nx4), .D (
         nx28447z1), .R (reset_int)) ;
    FDRE \reg_data_out(30)  (.Q (data_out_1_0[30]), .C (clk_int), .CE (nx4), .D (
         nx37422z1), .R (reset_int)) ;
    FDRE \reg_data_out(32)  (.Q (data_out_1_0[32]), .C (clk_int), .CE (nx4), .D (
         nx39416z1), .R (reset_int)) ;
    FDRE \reg_data_out(20)  (.Q (data_out_1_0[20]), .C (clk_int), .CE (nx4), .D (
         nx26453z1), .R (reset_int)) ;
    FDRE \reg_data_out(18)  (.Q (data_out_1_0[18]), .C (clk_int), .CE (nx4), .D (
         nx23460z1), .R (reset_int)) ;
    FDRE \reg_data_out(56)  (.Q (data_out_1_0[56]), .C (clk_int), .CE (nx4), .D (
         nx65342z1), .R (reset_int)) ;
    FDRE \reg_data_out(28)  (.Q (data_out_1_0[28]), .C (clk_int), .CE (nx4), .D (
         nx34429z1), .R (reset_int)) ;
    FDRE \reg_data_out(42)  (.Q (data_out_1_0[42]), .C (clk_int), .CE (nx4), .D (
         nx50385z1), .R (reset_int)) ;
    FDRE \reg_data_out(54)  (.Q (data_out_1_0[54]), .C (clk_int), .CE (nx4), .D (
         nx63348z1), .R (reset_int)) ;
    FDRE \reg_data_out(38)  (.Q (data_out_1_0[38]), .C (clk_int), .CE (nx4), .D (
         nx45398z1), .R (reset_int)) ;
    FDRE \reg_data_out(16)  (.Q (data_out_1_0[16]), .C (clk_int), .CE (nx4), .D (
         nx21466z1), .R (reset_int)) ;
    FDRE \reg_data_out(52)  (.Q (data_out_1_0[52]), .C (clk_int), .CE (nx4), .D (
         nx61354z1), .R (reset_int)) ;
    FDRE \reg_data_out(34)  (.Q (data_out_1_0[34]), .C (clk_int), .CE (nx4), .D (
         nx41410z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(63)  (.Q (data_out_1_0[63]), .C (
         clk_int), .CE (nx4), .D (nx63706z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(61)  (.Q (data_out_1_0[61]), .C (
         clk_int), .CE (nx4), .D (nx164z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(59)  (.Q (data_out_1_0[59]), .C (
         clk_int), .CE (nx4), .D (nx3157z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(57)  (.Q (data_out_1_0[57]), .C (
         clk_int), .CE (nx4), .D (nx5151z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(55)  (.Q (data_out_1_0[55]), .C (
         clk_int), .CE (nx4), .D (nx7145z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(53)  (.Q (data_out_1_0[53]), .C (
         clk_int), .CE (nx4), .D (nx9139z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(51)  (.Q (data_out_1_0[51]), .C (
         clk_int), .CE (nx4), .D (nx11133z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(49)  (.Q (data_out_1_0[49]), .C (
         clk_int), .CE (nx4), .D (nx14126z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(47)  (.Q (data_out_1_0[47]), .C (
         clk_int), .CE (nx4), .D (nx16120z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(45)  (.Q (data_out_1_0[45]), .C (
         clk_int), .CE (nx4), .D (nx18114z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(43)  (.Q (data_out_1_0[43]), .C (
         clk_int), .CE (nx4), .D (nx20108z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(41)  (.Q (data_out_1_0[41]), .C (
         clk_int), .CE (nx4), .D (nx22102z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(39)  (.Q (data_out_1_0[39]), .C (
         clk_int), .CE (nx4), .D (nx25095z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(37)  (.Q (data_out_1_0[37]), .C (
         clk_int), .CE (nx4), .D (nx27089z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(35)  (.Q (data_out_1_0[35]), .C (
         clk_int), .CE (nx4), .D (nx29083z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(33)  (.Q (data_out_1_0[33]), .C (
         clk_int), .CE (nx4), .D (nx31077z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(31)  (.Q (data_out_1_0[31]), .C (
         clk_int), .CE (nx4), .D (nx33071z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(29)  (.Q (data_out_1_0[29]), .C (
         clk_int), .CE (nx4), .D (nx36064z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(27)  (.Q (data_out_1_0[27]), .C (
         clk_int), .CE (nx4), .D (nx38058z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(25)  (.Q (data_out_1_0[25]), .C (
         clk_int), .CE (nx4), .D (nx40052z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(23)  (.Q (data_out_1_0[23]), .C (
         clk_int), .CE (nx4), .D (nx42046z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(21)  (.Q (data_out_1_0[21]), .C (
         clk_int), .CE (nx4), .D (nx44040z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(19)  (.Q (data_out_1_0[19]), .C (
         clk_int), .CE (nx4), .D (nx47033z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(17)  (.Q (data_out_1_0[17]), .C (
         clk_int), .CE (nx4), .D (nx49027z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(15)  (.Q (data_out_1_0[15]), .C (
         clk_int), .CE (nx4), .D (nx51021z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(13)  (.Q (data_out_1_0[13]), .C (
         clk_int), .CE (nx4), .D (nx53015z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(11)  (.Q (data_out_1_0[11]), .C (
         clk_int), .CE (nx4), .D (nx55009z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(9)  (.Q (data_out_1_0[9]), .C (clk_int)
         , .CE (nx4), .D (nx65314z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(7)  (.Q (data_out_1_0[7]), .C (clk_int)
         , .CE (nx4), .D (nx1772z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(5)  (.Q (data_out_1_0[5]), .C (clk_int)
         , .CE (nx4), .D (nx3766z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(3)  (.Q (data_out_1_0[3]), .C (clk_int)
         , .CE (nx4), .D (nx5760z1), .R (reset_int)) ;
    FDRE \i_output_tegister_reg_data_out(1)  (.Q (data_out_1_0[1]), .C (clk_int)
         , .CE (nx4), .D (nx7754z1), .R (reset_int)) ;
endmodule


module input_register_1 ( \p_plaintext(5)  , px3923, px3872, \p_plaintext(63)  , 
                          px3870, px3745, \p_plaintext(37)  , px3744, px3781, 
                          \p_plaintext(39)  , px3697, px3089, px3076, px3059, 
                          px3056, px3635, px3636, px3053, px3040, px3034, px3021, 
                          px3016, px3752, px3761, px3015, px3726, px3737, px3008, 
                          px3005, px3739, px3750, px2999, px2996, px2986, px2984, 
                          px2981, px3460, px3705, px3714, px2972, px2969, px2966, 
                          px3638, px3639, px2963, px3483, px3674, px3675, px2959, 
                          px2952, px2944, px2942, px2940, px3448, px3688, px3689, 
                          px2939, px3716, px3717, px2935, px3626, px3627, px2934, 
                          px3623, px3624, px2933, px2928, px2926, px3702, px3703, 
                          px2925, px3657, px3658, px2924, px3665, px3666, px2921, 
                          px2913, px2912, px2908, px2906, px2898, px3584, px3585, 
                          px2897, px3335, px3590, px3591, px2896, px2894, px2892, 
                          px2890, px3649, px3650, px2887, px3632, px3647, px2886, 
                          px2884, px3338, px3546, px3547, px2879, px3408, px3652, 
                          px3667, px2878, px3615, px3630, px2877, px3543, px3544, 
                          px2872, px2870, px3405, px3406, px2867, px3523, px3534, 
                          px2866, px3596, px3607, px2865, px3587, px3588, px2860, 
                          px3559, px3560, px2859, px3562, px3563, px2858, px3514, 
                          px3515, px2847, px3511, px3512, px2846, px3359, px3565, 
                          px3576, px2845, px3724, px3886, px2844, px3582, px3611, 
                          px2841, px2835, px3392, px3403, px2827, px2823, px2821, 
                          px3436, px3437, px2812, px2810, px3442, px3443, px2803, 
                          px2801, px3421, px3422, px2797, px3506, px3521, px2796, 
                          px2794, px3536, px3551, px2793, px3439, px3440, px2780, 
                          px3454, px3455, px2777, px3433, px3434, px2773, px2765, 
                          px3504, px3723, px2764, px3451, px3452, px2763, px3410, 
                          px3411, px2760, px2751, px3315, px3316, px2741, px3321, 
                          px3322, px2733, px2731, px3304, px3305, px2729, px3332, 
                          px3333, px2723, px2719, px3425, px3444, px2712, px3341, 
                          px3342, px2711, px2709, px2706, px3373, px3374, px2703, 
                          px3353, px3354, px2702, px3307, px3308, px2698, px2694, 
                          px2732, px2881, px3090, px3313, px3328, px2683, px2766, 
                          px2927, px3136, px3330, px3349, px2682, px2680, px2678, 
                          px2672, px2670, px2710, px2871, px3077, px3283, px3294, 
                          px2669, px2720, px2893, px3060, px3296, px3311, px2668, 
                          px2664, px2658, px2656, px2654, px2646, px2644, px2671, 
                          px2855, px3010, px3216, px3217, px2643, px3206, px3207, 
                          px2642, px2640, px2638, px2647, px2832, px3054, px3197, 
                          px3198, px2637, px3191, px3192, px2634, px2630, px2628, 
                          px2659, px2824, px2982, px3235, px3236, px2623, px2695, 
                          px2798, px2997, px3278, px3279, px2622, px2681, px2795, 
                          px2987, px3261, px3262, px2621, px2665, px2820, px2973, 
                          px3232, px3233, px2618, px2615, px2613, px2611, px2657, 
                          px2822, px2967, px3226, px3227, px2608, px2655, px2818, 
                          px2970, px3229, px3230, px2607, px2639, px2807, px3022, 
                          px3172, px3173, px2606, px3183, px3184, px2605, px2601, 
                          px2593, px2591, px2587, px2585, px2641, px2828, px2953, 
                          px3187, px3202, px2582, px2707, px2868, px3057, px3221, 
                          px3222, px2579, px2575, px2573, px2592, px2786, px2945, 
                          px3160, px3161, px2570, px2679, px2790, px2985, px3245, 
                          px3280, px2569, px2629, px2802, px3017, px3170, px3185, 
                          px2566, px2594, px2772, px2929, px3138, px3149, px2563, 
                          px2588, px2768, px2941, px3151, px3152, px2558, px2586, 
                          px2770, px2943, px3154, px3155, px2557, px2555, px2551, 
                          px2602, px2748, px2914, px3119, px3120, px2538, px2574, 
                          px2734, px2885, px3095, px3096, px2537, px2576, px2742, 
                          px2891, px3092, px3093, px2534, px2708, px2869, px3058, 
                          px3281, px3503, px2533, px2552, px2728, px2895, px3073, 
                          px3074, px2528, px2612, px2746, px2907, px3109, px3110, 
                          px2523, px2556, px2730, px2899, px3068, px3069, px2522, 
                          px2614, px2752, px2909, px3112, px3113, px2521, px2520, 
                          px2673, px2857, px3006, px3007, px2514, px2508, px2645, 
                          px2836, px3035, px3036, px2507, px2498, px2631, px2811, 
                          px3041, px3052, px2497, p_nbus_key_in_int, 
                          \p_key_samp(1)  , \p_key_samp(2)  , \p_key_samp(3)  , 
                          \p_key_samp(4)  , \p_key_samp(5)  , \p_key_samp(6)  , 
                          \p_key_samp(7)  , \p_key_samp(9)  , \p_key_samp(10)  , 
                          \p_key_samp(11)  , \p_key_samp(12)  , \p_key_samp(13)  , 
                          \p_key_samp(14)  , \p_key_samp(15)  , \p_key_samp(17)  , 
                          \p_key_samp(18)  , \p_key_samp(19)  , \p_key_samp(20)  , 
                          \p_key_samp(21)  , \p_key_samp(22)  , \p_key_samp(23)  , 
                          \p_key_samp(25)  , \p_key_samp(26)  , \p_key_samp(27)  , 
                          \p_key_samp(28)  , \p_key_samp(29)  , \p_key_samp(30)  , 
                          \p_key_samp(31)  , \p_key_samp(33)  , \p_key_samp(34)  , 
                          \p_key_samp(35)  , \p_key_samp(36)  , \p_key_samp(37)  , 
                          \p_key_samp(38)  , \p_key_samp(39)  , \p_key_samp(41)  , 
                          \p_key_samp(42)  , \p_key_samp(43)  , \p_key_samp(44)  , 
                          \p_key_samp(45)  , \p_key_samp(46)  , \p_key_samp(47)  , 
                          \p_key_samp(49)  , \p_key_samp(50)  , \p_key_samp(51)  , 
                          \p_key_samp(52)  , \p_key_samp(53)  , \p_key_samp(54)  , 
                          \p_key_samp(55)  , \p_key_samp(57)  , \p_key_samp(58)  , 
                          \p_key_samp(59)  , \p_key_samp(60)  , \p_key_samp(61)  , 
                          \p_key_samp(62)  , p_reset_int, p_load_int, p_clk_int, 
                          \p_key_samp(63)   ) ;

    input \p_plaintext(5)   ;
    output px3923 ;
    output px3872 ;
    input \p_plaintext(63)   ;
    output px3870 ;
    input px3745 ;
    input \p_plaintext(37)   ;
    output px3744 ;
    input px3781 ;
    input \p_plaintext(39)   ;
    output px3697 ;
    output px3089 ;
    output px3076 ;
    output px3059 ;
    output px3056 ;
    input px3635 ;
    input px3636 ;
    output px3053 ;
    output px3040 ;
    output px3034 ;
    output px3021 ;
    output px3016 ;
    input px3752 ;
    input px3761 ;
    output px3015 ;
    input px3726 ;
    input px3737 ;
    output px3008 ;
    output px3005 ;
    input px3739 ;
    input px3750 ;
    output px2999 ;
    output px2996 ;
    output px2986 ;
    output px2984 ;
    output px2981 ;
    input px3460 ;
    input px3705 ;
    input px3714 ;
    output px2972 ;
    output px2969 ;
    output px2966 ;
    input px3638 ;
    input px3639 ;
    output px2963 ;
    input px3483 ;
    input px3674 ;
    input px3675 ;
    output px2959 ;
    output px2952 ;
    output px2944 ;
    output px2942 ;
    output px2940 ;
    input px3448 ;
    input px3688 ;
    input px3689 ;
    output px2939 ;
    input px3716 ;
    input px3717 ;
    output px2935 ;
    input px3626 ;
    input px3627 ;
    output px2934 ;
    input px3623 ;
    input px3624 ;
    output px2933 ;
    output px2928 ;
    output px2926 ;
    input px3702 ;
    input px3703 ;
    output px2925 ;
    input px3657 ;
    input px3658 ;
    output px2924 ;
    input px3665 ;
    input px3666 ;
    output px2921 ;
    output px2913 ;
    output px2912 ;
    output px2908 ;
    output px2906 ;
    output px2898 ;
    input px3584 ;
    input px3585 ;
    output px2897 ;
    input px3335 ;
    input px3590 ;
    input px3591 ;
    output px2896 ;
    output px2894 ;
    output px2892 ;
    output px2890 ;
    input px3649 ;
    input px3650 ;
    output px2887 ;
    input px3632 ;
    input px3647 ;
    output px2886 ;
    output px2884 ;
    input px3338 ;
    input px3546 ;
    input px3547 ;
    output px2879 ;
    input px3408 ;
    input px3652 ;
    input px3667 ;
    output px2878 ;
    input px3615 ;
    input px3630 ;
    output px2877 ;
    input px3543 ;
    input px3544 ;
    output px2872 ;
    output px2870 ;
    input px3405 ;
    input px3406 ;
    output px2867 ;
    input px3523 ;
    input px3534 ;
    output px2866 ;
    input px3596 ;
    input px3607 ;
    output px2865 ;
    input px3587 ;
    input px3588 ;
    output px2860 ;
    input px3559 ;
    input px3560 ;
    output px2859 ;
    input px3562 ;
    input px3563 ;
    output px2858 ;
    input px3514 ;
    input px3515 ;
    output px2847 ;
    input px3511 ;
    input px3512 ;
    output px2846 ;
    input px3359 ;
    input px3565 ;
    input px3576 ;
    output px2845 ;
    input px3724 ;
    input px3886 ;
    output px2844 ;
    input px3582 ;
    input px3611 ;
    output px2841 ;
    output px2835 ;
    input px3392 ;
    input px3403 ;
    output px2827 ;
    output px2823 ;
    output px2821 ;
    input px3436 ;
    input px3437 ;
    output px2812 ;
    output px2810 ;
    input px3442 ;
    input px3443 ;
    output px2803 ;
    output px2801 ;
    input px3421 ;
    input px3422 ;
    output px2797 ;
    input px3506 ;
    input px3521 ;
    output px2796 ;
    output px2794 ;
    input px3536 ;
    input px3551 ;
    output px2793 ;
    input px3439 ;
    input px3440 ;
    output px2780 ;
    input px3454 ;
    input px3455 ;
    output px2777 ;
    input px3433 ;
    input px3434 ;
    output px2773 ;
    output px2765 ;
    input px3504 ;
    input px3723 ;
    output px2764 ;
    input px3451 ;
    input px3452 ;
    output px2763 ;
    input px3410 ;
    input px3411 ;
    output px2760 ;
    output px2751 ;
    input px3315 ;
    input px3316 ;
    output px2741 ;
    input px3321 ;
    input px3322 ;
    output px2733 ;
    output px2731 ;
    input px3304 ;
    input px3305 ;
    output px2729 ;
    input px3332 ;
    input px3333 ;
    output px2723 ;
    output px2719 ;
    input px3425 ;
    input px3444 ;
    output px2712 ;
    input px3341 ;
    input px3342 ;
    output px2711 ;
    output px2709 ;
    output px2706 ;
    input px3373 ;
    input px3374 ;
    output px2703 ;
    input px3353 ;
    input px3354 ;
    output px2702 ;
    input px3307 ;
    input px3308 ;
    output px2698 ;
    output px2694 ;
    input px2732 ;
    input px2881 ;
    input px3090 ;
    input px3313 ;
    input px3328 ;
    output px2683 ;
    input px2766 ;
    input px2927 ;
    input px3136 ;
    input px3330 ;
    input px3349 ;
    output px2682 ;
    output px2680 ;
    output px2678 ;
    output px2672 ;
    output px2670 ;
    input px2710 ;
    input px2871 ;
    input px3077 ;
    input px3283 ;
    input px3294 ;
    output px2669 ;
    input px2720 ;
    input px2893 ;
    input px3060 ;
    input px3296 ;
    input px3311 ;
    output px2668 ;
    output px2664 ;
    output px2658 ;
    output px2656 ;
    output px2654 ;
    output px2646 ;
    output px2644 ;
    input px2671 ;
    input px2855 ;
    input px3010 ;
    input px3216 ;
    input px3217 ;
    output px2643 ;
    input px3206 ;
    input px3207 ;
    output px2642 ;
    output px2640 ;
    output px2638 ;
    input px2647 ;
    input px2832 ;
    input px3054 ;
    input px3197 ;
    input px3198 ;
    output px2637 ;
    input px3191 ;
    input px3192 ;
    output px2634 ;
    output px2630 ;
    output px2628 ;
    input px2659 ;
    input px2824 ;
    input px2982 ;
    input px3235 ;
    input px3236 ;
    output px2623 ;
    input px2695 ;
    input px2798 ;
    input px2997 ;
    input px3278 ;
    input px3279 ;
    output px2622 ;
    input px2681 ;
    input px2795 ;
    input px2987 ;
    input px3261 ;
    input px3262 ;
    output px2621 ;
    input px2665 ;
    input px2820 ;
    input px2973 ;
    input px3232 ;
    input px3233 ;
    output px2618 ;
    output px2615 ;
    output px2613 ;
    output px2611 ;
    input px2657 ;
    input px2822 ;
    input px2967 ;
    input px3226 ;
    input px3227 ;
    output px2608 ;
    input px2655 ;
    input px2818 ;
    input px2970 ;
    input px3229 ;
    input px3230 ;
    output px2607 ;
    input px2639 ;
    input px2807 ;
    input px3022 ;
    input px3172 ;
    input px3173 ;
    output px2606 ;
    input px3183 ;
    input px3184 ;
    output px2605 ;
    output px2601 ;
    output px2593 ;
    output px2591 ;
    output px2587 ;
    output px2585 ;
    input px2641 ;
    input px2828 ;
    input px2953 ;
    input px3187 ;
    input px3202 ;
    output px2582 ;
    input px2707 ;
    input px2868 ;
    input px3057 ;
    input px3221 ;
    input px3222 ;
    output px2579 ;
    output px2575 ;
    output px2573 ;
    input px2592 ;
    input px2786 ;
    input px2945 ;
    input px3160 ;
    input px3161 ;
    output px2570 ;
    input px2679 ;
    input px2790 ;
    input px2985 ;
    input px3245 ;
    input px3280 ;
    output px2569 ;
    input px2629 ;
    input px2802 ;
    input px3017 ;
    input px3170 ;
    input px3185 ;
    output px2566 ;
    input px2594 ;
    input px2772 ;
    input px2929 ;
    input px3138 ;
    input px3149 ;
    output px2563 ;
    input px2588 ;
    input px2768 ;
    input px2941 ;
    input px3151 ;
    input px3152 ;
    output px2558 ;
    input px2586 ;
    input px2770 ;
    input px2943 ;
    input px3154 ;
    input px3155 ;
    output px2557 ;
    output px2555 ;
    output px2551 ;
    input px2602 ;
    input px2748 ;
    input px2914 ;
    input px3119 ;
    input px3120 ;
    output px2538 ;
    input px2574 ;
    input px2734 ;
    input px2885 ;
    input px3095 ;
    input px3096 ;
    output px2537 ;
    input px2576 ;
    input px2742 ;
    input px2891 ;
    input px3092 ;
    input px3093 ;
    output px2534 ;
    input px2708 ;
    input px2869 ;
    input px3058 ;
    input px3281 ;
    input px3503 ;
    output px2533 ;
    input px2552 ;
    input px2728 ;
    input px2895 ;
    input px3073 ;
    input px3074 ;
    output px2528 ;
    input px2612 ;
    input px2746 ;
    input px2907 ;
    input px3109 ;
    input px3110 ;
    output px2523 ;
    input px2556 ;
    input px2730 ;
    input px2899 ;
    input px3068 ;
    input px3069 ;
    output px2522 ;
    input px2614 ;
    input px2752 ;
    input px2909 ;
    input px3112 ;
    input px3113 ;
    output px2521 ;
    input px2520 ;
    input px2673 ;
    input px2857 ;
    input px3006 ;
    input px3007 ;
    output px2514 ;
    input px2508 ;
    input px2645 ;
    input px2836 ;
    input px3035 ;
    input px3036 ;
    output px2507 ;
    input px2498 ;
    input px2631 ;
    input px2811 ;
    input px3041 ;
    input px3052 ;
    output px2497 ;
    input [63:8]p_nbus_key_in_int ;
    output \p_key_samp(1)   ;
    output \p_key_samp(2)   ;
    output \p_key_samp(3)   ;
    output \p_key_samp(4)   ;
    output \p_key_samp(5)   ;
    output \p_key_samp(6)   ;
    output \p_key_samp(7)   ;
    output \p_key_samp(9)   ;
    output \p_key_samp(10)   ;
    output \p_key_samp(11)   ;
    output \p_key_samp(12)   ;
    output \p_key_samp(13)   ;
    output \p_key_samp(14)   ;
    output \p_key_samp(15)   ;
    output \p_key_samp(17)   ;
    output \p_key_samp(18)   ;
    output \p_key_samp(19)   ;
    output \p_key_samp(20)   ;
    output \p_key_samp(21)   ;
    output \p_key_samp(22)   ;
    output \p_key_samp(23)   ;
    output \p_key_samp(25)   ;
    output \p_key_samp(26)   ;
    output \p_key_samp(27)   ;
    output \p_key_samp(28)   ;
    output \p_key_samp(29)   ;
    output \p_key_samp(30)   ;
    output \p_key_samp(31)   ;
    output \p_key_samp(33)   ;
    output \p_key_samp(34)   ;
    output \p_key_samp(35)   ;
    output \p_key_samp(36)   ;
    output \p_key_samp(37)   ;
    output \p_key_samp(38)   ;
    output \p_key_samp(39)   ;
    output \p_key_samp(41)   ;
    output \p_key_samp(42)   ;
    output \p_key_samp(43)   ;
    output \p_key_samp(44)   ;
    output \p_key_samp(45)   ;
    output \p_key_samp(46)   ;
    output \p_key_samp(47)   ;
    output \p_key_samp(49)   ;
    output \p_key_samp(50)   ;
    output \p_key_samp(51)   ;
    output \p_key_samp(52)   ;
    output \p_key_samp(53)   ;
    output \p_key_samp(54)   ;
    output \p_key_samp(55)   ;
    output \p_key_samp(57)   ;
    output \p_key_samp(58)   ;
    output \p_key_samp(59)   ;
    output \p_key_samp(60)   ;
    output \p_key_samp(61)   ;
    output \p_key_samp(62)   ;
    input p_reset_int ;
    input p_load_int ;
    input p_clk_int ;
    output \p_key_samp(63)   ;




    FDRE \reg_data_out(63)  (.Q (\p_key_samp(63)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[8]), .R (p_reset_int)) ;
    FDRE \reg_data_out(62)  (.Q (\p_key_samp(62)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[9]), .R (p_reset_int)) ;
    FDRE \reg_data_out(61)  (.Q (\p_key_samp(61)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[10]), .R (p_reset_int)) ;
    FDRE \reg_data_out(60)  (.Q (\p_key_samp(60)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[11]), .R (p_reset_int)) ;
    FDRE \reg_data_out(59)  (.Q (\p_key_samp(59)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[12]), .R (p_reset_int)) ;
    FDRE \reg_data_out(58)  (.Q (\p_key_samp(58)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[13]), .R (p_reset_int)) ;
    FDRE \reg_data_out(57)  (.Q (\p_key_samp(57)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[14]), .R (p_reset_int)) ;
    FDRE \reg_data_out(55)  (.Q (\p_key_samp(55)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[15]), .R (p_reset_int)) ;
    FDRE \reg_data_out(54)  (.Q (\p_key_samp(54)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[16]), .R (p_reset_int)) ;
    FDRE \reg_data_out(53)  (.Q (\p_key_samp(53)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[17]), .R (p_reset_int)) ;
    FDRE \reg_data_out(52)  (.Q (\p_key_samp(52)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[18]), .R (p_reset_int)) ;
    FDRE \reg_data_out(51)  (.Q (\p_key_samp(51)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[19]), .R (p_reset_int)) ;
    FDRE \reg_data_out(50)  (.Q (\p_key_samp(50)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[20]), .R (p_reset_int)) ;
    FDRE \reg_data_out(49)  (.Q (\p_key_samp(49)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[21]), .R (p_reset_int)) ;
    FDRE \reg_data_out(47)  (.Q (\p_key_samp(47)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[22]), .R (p_reset_int)) ;
    FDRE \reg_data_out(46)  (.Q (\p_key_samp(46)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[23]), .R (p_reset_int)) ;
    FDRE \reg_data_out(45)  (.Q (\p_key_samp(45)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[24]), .R (p_reset_int)) ;
    FDRE \reg_data_out(44)  (.Q (\p_key_samp(44)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[25]), .R (p_reset_int)) ;
    FDRE \reg_data_out(43)  (.Q (\p_key_samp(43)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[26]), .R (p_reset_int)) ;
    FDRE \reg_data_out(42)  (.Q (\p_key_samp(42)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[27]), .R (p_reset_int)) ;
    FDRE \reg_data_out(41)  (.Q (\p_key_samp(41)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[28]), .R (p_reset_int)) ;
    FDRE \reg_data_out(39)  (.Q (\p_key_samp(39)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[29]), .R (p_reset_int)) ;
    FDRE \reg_data_out(38)  (.Q (\p_key_samp(38)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[30]), .R (p_reset_int)) ;
    FDRE \reg_data_out(37)  (.Q (\p_key_samp(37)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[31]), .R (p_reset_int)) ;
    FDRE \reg_data_out(36)  (.Q (\p_key_samp(36)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[32]), .R (p_reset_int)) ;
    FDRE \reg_data_out(35)  (.Q (\p_key_samp(35)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[33]), .R (p_reset_int)) ;
    FDRE \reg_data_out(34)  (.Q (\p_key_samp(34)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[34]), .R (p_reset_int)) ;
    FDRE \reg_data_out(33)  (.Q (\p_key_samp(33)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[35]), .R (p_reset_int)) ;
    FDRE \reg_data_out(31)  (.Q (\p_key_samp(31)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[36]), .R (p_reset_int)) ;
    FDRE \reg_data_out(30)  (.Q (\p_key_samp(30)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[37]), .R (p_reset_int)) ;
    FDRE \reg_data_out(29)  (.Q (\p_key_samp(29)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[38]), .R (p_reset_int)) ;
    FDRE \reg_data_out(28)  (.Q (\p_key_samp(28)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[39]), .R (p_reset_int)) ;
    FDRE \reg_data_out(27)  (.Q (\p_key_samp(27)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[40]), .R (p_reset_int)) ;
    FDRE \reg_data_out(26)  (.Q (\p_key_samp(26)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[41]), .R (p_reset_int)) ;
    FDRE \reg_data_out(25)  (.Q (\p_key_samp(25)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[42]), .R (p_reset_int)) ;
    FDRE \reg_data_out(23)  (.Q (\p_key_samp(23)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[43]), .R (p_reset_int)) ;
    FDRE \reg_data_out(22)  (.Q (\p_key_samp(22)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[44]), .R (p_reset_int)) ;
    FDRE \reg_data_out(21)  (.Q (\p_key_samp(21)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[45]), .R (p_reset_int)) ;
    FDRE \reg_data_out(20)  (.Q (\p_key_samp(20)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[46]), .R (p_reset_int)) ;
    FDRE \reg_data_out(19)  (.Q (\p_key_samp(19)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[47]), .R (p_reset_int)) ;
    FDRE \reg_data_out(18)  (.Q (\p_key_samp(18)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[48]), .R (p_reset_int)) ;
    FDRE \reg_data_out(17)  (.Q (\p_key_samp(17)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[49]), .R (p_reset_int)) ;
    FDRE \reg_data_out(15)  (.Q (\p_key_samp(15)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[50]), .R (p_reset_int)) ;
    FDRE \reg_data_out(14)  (.Q (\p_key_samp(14)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[51]), .R (p_reset_int)) ;
    FDRE \reg_data_out(13)  (.Q (\p_key_samp(13)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[52]), .R (p_reset_int)) ;
    FDRE \reg_data_out(12)  (.Q (\p_key_samp(12)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[53]), .R (p_reset_int)) ;
    FDRE \reg_data_out(11)  (.Q (\p_key_samp(11)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[54]), .R (p_reset_int)) ;
    FDRE \reg_data_out(10)  (.Q (\p_key_samp(10)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[55]), .R (p_reset_int)) ;
    FDRE \reg_data_out(9)  (.Q (\p_key_samp(9)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[56]), .R (p_reset_int)) ;
    FDRE \reg_data_out(7)  (.Q (\p_key_samp(7)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[57]), .R (p_reset_int)) ;
    FDRE \reg_data_out(6)  (.Q (\p_key_samp(6)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[58]), .R (p_reset_int)) ;
    FDRE \reg_data_out(5)  (.Q (\p_key_samp(5)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[59]), .R (p_reset_int)) ;
    FDRE \reg_data_out(4)  (.Q (\p_key_samp(4)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[60]), .R (p_reset_int)) ;
    FDRE \reg_data_out(3)  (.Q (\p_key_samp(3)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[61]), .R (p_reset_int)) ;
    FDRE \reg_data_out(2)  (.Q (\p_key_samp(2)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[62]), .R (p_reset_int)) ;
    FDRE \reg_data_out(1)  (.Q (\p_key_samp(1)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_key_in_int[63]), .R (p_reset_int)) ;
    LUT6 ix36838z39819 (.O (px2497), .I0 (\p_key_samp(15)  ), .I1 (px3052), .I2 (
         px3041), .I3 (px2811), .I4 (px2631), .I5 (px2498)) ;
         defparam ix36838z39819.INIT = 64'h9669699669969669;
    LUT6 ix34842z28344 (.O (px2507), .I0 (\p_key_samp(12)  ), .I1 (px3036), .I2 (
         px3035), .I3 (px2836), .I4 (px2645), .I5 (px2508)) ;
         defparam ix34842z28344.INIT = 64'h6996966996696996;
    LUT6 ix33848z28344 (.O (px2514), .I0 (\p_key_samp(21)  ), .I1 (px3007), .I2 (
         px3006), .I3 (px2857), .I4 (px2673), .I5 (px2520)) ;
         defparam ix33848z28344.INIT = 64'h6996966996696996;
    LUT6 ix32854z39819 (.O (px2521), .I0 (\p_key_samp(28)  ), .I1 (px3113), .I2 (
         px3112), .I3 (px2909), .I4 (px2752), .I5 (px2614)) ;
         defparam ix32854z39819.INIT = 64'h9669699669969669;
    LUT6 ix32853z39819 (.O (px2522), .I0 (\p_key_samp(62)  ), .I1 (px3069), .I2 (
         px3068), .I3 (px2899), .I4 (px2730), .I5 (px2556)) ;
         defparam ix32853z39819.INIT = 64'h9669699669969669;
    LUT6 ix32852z28344 (.O (px2523), .I0 (\p_key_samp(31)  ), .I1 (px3110), .I2 (
         px3109), .I3 (px2907), .I4 (px2746), .I5 (px2612)) ;
         defparam ix32852z28344.INIT = 64'h6996966996696996;
    LUT6 ix32847z39819 (.O (px2528), .I0 (\p_key_samp(38)  ), .I1 (px3074), .I2 (
         px3073), .I3 (px2895), .I4 (px2728), .I5 (px2552)) ;
         defparam ix32847z39819.INIT = 64'h9669699669969669;
    LUT6 ix31855z39819 (.O (px2533), .I0 (\p_key_samp(13)  ), .I1 (px3503), .I2 (
         px3281), .I3 (px3058), .I4 (px2869), .I5 (px2708)) ;
         defparam ix31855z39819.INIT = 64'h9669699669969669;
    LUT6 ix31854z28344 (.O (px2534), .I0 (\p_key_samp(55)  ), .I1 (px3093), .I2 (
         px3092), .I3 (px2891), .I4 (px2742), .I5 (px2576)) ;
         defparam ix31854z28344.INIT = 64'h6996966996696996;
    LUT6 ix31851z39819 (.O (px2537), .I0 (\p_key_samp(4)  ), .I1 (px3096), .I2 (
         px3095), .I3 (px2885), .I4 (px2734), .I5 (px2574)) ;
         defparam ix31851z39819.INIT = 64'h9669699669969669;
    LUT6 ix31850z39819 (.O (px2538), .I0 (\p_key_samp(45)  ), .I1 (px3120), .I2 (
         px3119), .I3 (px2914), .I4 (px2748), .I5 (px2602)) ;
         defparam ix31850z39819.INIT = 64'h9669699669969669;
    LUT6 ix29863z39819 (.O (px2551), .I0 (\p_key_samp(60)  ), .I1 (px3074), .I2 (
         px3073), .I3 (px2895), .I4 (px2728), .I5 (px2552)) ;
         defparam ix29863z39819.INIT = 64'h9669699669969669;
    LUT6 ix29859z39819 (.O (px2555), .I0 (\p_key_samp(17)  ), .I1 (px3069), .I2 (
         px3068), .I3 (px2899), .I4 (px2730), .I5 (px2556)) ;
         defparam ix29859z39819.INIT = 64'h9669699669969669;
    LUT6 ix29857z28344 (.O (px2557), .I0 (\p_key_samp(34)  ), .I1 (px3155), .I2 (
         px3154), .I3 (px2943), .I4 (px2770), .I5 (px2586)) ;
         defparam ix29857z28344.INIT = 64'h6996966996696996;
    LUT6 ix29856z28344 (.O (px2558), .I0 (\p_key_samp(3)  ), .I1 (px3152), .I2 (
         px3151), .I3 (px2941), .I4 (px2768), .I5 (px2588)) ;
         defparam ix29856z28344.INIT = 64'h6996966996696996;
    LUT6 ix28864z28344 (.O (px2563), .I0 (\p_key_samp(19)  ), .I1 (px3149), .I2 (
         px3138), .I3 (px2929), .I4 (px2772), .I5 (px2594)) ;
         defparam ix28864z28344.INIT = 64'h6996966996696996;
    LUT6 ix28861z39819 (.O (px2566), .I0 (\p_key_samp(1)  ), .I1 (px3185), .I2 (
         px3170), .I3 (px3017), .I4 (px2802), .I5 (px2629)) ;
         defparam ix28861z39819.INIT = 64'h9669699669969669;
    LUT6 ix28858z39819 (.O (px2569), .I0 (\p_key_samp(18)  ), .I1 (px3280), .I2 (
         px3245), .I3 (px2985), .I4 (px2790), .I5 (px2679)) ;
         defparam ix28858z39819.INIT = 64'h9669699669969669;
    LUT6 ix27870z39819 (.O (px2570), .I0 (\p_key_samp(25)  ), .I1 (px3161), .I2 (
         px3160), .I3 (px2945), .I4 (px2786), .I5 (px2592)) ;
         defparam ix27870z39819.INIT = 64'h9669699669969669;
    LUT6 ix27867z39819 (.O (px2573), .I0 (\p_key_samp(54)  ), .I1 (px3096), .I2 (
         px3095), .I3 (px2885), .I4 (px2734), .I5 (px2574)) ;
         defparam ix27867z39819.INIT = 64'h9669699669969669;
    LUT6 ix27865z28344 (.O (px2575), .I0 (\p_key_samp(47)  ), .I1 (px3093), .I2 (
         px3092), .I3 (px2891), .I4 (px2742), .I5 (px2576)) ;
         defparam ix27865z28344.INIT = 64'h6996966996696996;
    LUT6 ix27861z39819 (.O (px2579), .I0 (\p_key_samp(7)  ), .I1 (px3222), .I2 (
         px3221), .I3 (px3057), .I4 (px2868), .I5 (px2707)) ;
         defparam ix27861z39819.INIT = 64'h9669699669969669;
    LUT6 ix26871z39819 (.O (px2582), .I0 (\p_key_samp(30)  ), .I1 (px3202), .I2 (
         px3187), .I3 (px2953), .I4 (px2828), .I5 (px2641)) ;
         defparam ix26871z39819.INIT = 64'h9669699669969669;
    LUT6 ix26868z28344 (.O (px2585), .I0 (\p_key_samp(59)  ), .I1 (px3155), .I2 (
         px3154), .I3 (px2943), .I4 (px2770), .I5 (px2586)) ;
         defparam ix26868z28344.INIT = 64'h6996966996696996;
    LUT6 ix26866z28344 (.O (px2587), .I0 (\p_key_samp(33)  ), .I1 (px3152), .I2 (
         px3151), .I3 (px2941), .I4 (px2768), .I5 (px2588)) ;
         defparam ix26866z28344.INIT = 64'h6996966996696996;
    LUT6 ix25875z39819 (.O (px2591), .I0 (\p_key_samp(50)  ), .I1 (px3161), .I2 (
         px3160), .I3 (px2945), .I4 (px2786), .I5 (px2592)) ;
         defparam ix25875z39819.INIT = 64'h9669699669969669;
    LUT6 ix25873z28344 (.O (px2593), .I0 (\p_key_samp(27)  ), .I1 (px3149), .I2 (
         px3138), .I3 (px2929), .I4 (px2772), .I5 (px2594)) ;
         defparam ix25873z28344.INIT = 64'h6996966996696996;
    LUT6 ix23879z39819 (.O (px2601), .I0 (\p_key_samp(29)  ), .I1 (px3120), .I2 (
         px3119), .I3 (px2914), .I4 (px2748), .I5 (px2602)) ;
         defparam ix23879z39819.INIT = 64'h9669699669969669;
    LUT6 ix23875z39819 (.O (px2605), .I0 (\p_key_samp(35)  ), .I1 (px3184), .I2 (
         px3183), .I3 (px3041), .I4 (px2811), .I5 (px2631)) ;
         defparam ix23875z39819.INIT = 64'h9669699669969669;
    LUT6 ix23874z39819 (.O (px2606), .I0 (\p_key_samp(10)  ), .I1 (px3173), .I2 (
         px3172), .I3 (px3022), .I4 (px2807), .I5 (px2639)) ;
         defparam ix23874z39819.INIT = 64'h9669699669969669;
    LUT6 ix23873z39819 (.O (px2607), .I0 (\p_key_samp(59)  ), .I1 (px3230), .I2 (
         px3229), .I3 (px2970), .I4 (px2818), .I5 (px2655)) ;
         defparam ix23873z39819.INIT = 64'h9669699669969669;
    LUT6 ix23872z28344 (.O (px2608), .I0 (\p_key_samp(58)  ), .I1 (px3227), .I2 (
         px3226), .I3 (px2967), .I4 (px2822), .I5 (px2657)) ;
         defparam ix23872z28344.INIT = 64'h6996966996696996;
    LUT6 ix22882z28344 (.O (px2611), .I0 (\p_key_samp(20)  ), .I1 (px3110), .I2 (
         px3109), .I3 (px2907), .I4 (px2746), .I5 (px2612)) ;
         defparam ix22882z28344.INIT = 64'h6996966996696996;
    LUT6 ix22880z39819 (.O (px2613), .I0 (\p_key_samp(15)  ), .I1 (px3113), .I2 (
         px3112), .I3 (px2909), .I4 (px2752), .I5 (px2614)) ;
         defparam ix22880z39819.INIT = 64'h9669699669969669;
    LUT6 ix22878z39819 (.O (px2615), .I0 (\p_key_samp(6)  ), .I1 (px3503), .I2 (
         px3281), .I3 (px3058), .I4 (px2869), .I5 (px2708)) ;
         defparam ix22878z39819.INIT = 64'h9669699669969669;
    LUT6 ix22875z28344 (.O (px2618), .I0 (\p_key_samp(34)  ), .I1 (px3233), .I2 (
         px3232), .I3 (px2973), .I4 (px2820), .I5 (px2665)) ;
         defparam ix22875z28344.INIT = 64'h6996966996696996;
    LUT6 ix21885z39819 (.O (px2621), .I0 (\p_key_samp(17)  ), .I1 (px3262), .I2 (
         px3261), .I3 (px2987), .I4 (px2795), .I5 (px2681)) ;
         defparam ix21885z39819.INIT = 64'h9669699669969669;
    LUT6 ix21884z28344 (.O (px2622), .I0 (\p_key_samp(43)  ), .I1 (px3279), .I2 (
         px3278), .I3 (px2997), .I4 (px2798), .I5 (px2695)) ;
         defparam ix21884z28344.INIT = 64'h6996966996696996;
    LUT6 ix21883z39819 (.O (px2623), .I0 (\p_key_samp(11)  ), .I1 (px3236), .I2 (
         px3235), .I3 (px2982), .I4 (px2824), .I5 (px2659)) ;
         defparam ix21883z39819.INIT = 64'h9669699669969669;
    LUT6 ix21878z39819 (.O (px2628), .I0 (\p_key_samp(11)  ), .I1 (px3185), .I2 (
         px3170), .I3 (px3017), .I4 (px2802), .I5 (px2629)) ;
         defparam ix21878z39819.INIT = 64'h9669699669969669;
    LUT6 ix20889z39819 (.O (px2630), .I0 (\p_key_samp(20)  ), .I1 (px3184), .I2 (
         px3183), .I3 (px3041), .I4 (px2811), .I5 (px2631)) ;
         defparam ix20889z39819.INIT = 64'h9669699669969669;
    LUT6 ix20885z28344 (.O (px2634), .I0 (\p_key_samp(38)  ), .I1 (px3192), .I2 (
         px3191), .I3 (px3035), .I4 (px2836), .I5 (px2645)) ;
         defparam ix20885z28344.INIT = 64'h6996966996696996;
    LUT6 ix20882z39819 (.O (px2637), .I0 (\p_key_samp(31)  ), .I1 (px3198), .I2 (
         px3197), .I3 (px3054), .I4 (px2832), .I5 (px2647)) ;
         defparam ix20882z39819.INIT = 64'h9669699669969669;
    LUT6 ix20881z39819 (.O (px2638), .I0 (\p_key_samp(14)  ), .I1 (px3173), .I2 (
         px3172), .I3 (px3022), .I4 (px2807), .I5 (px2639)) ;
         defparam ix20881z39819.INIT = 64'h9669699669969669;
    LUT6 ix19892z39819 (.O (px2640), .I0 (\p_key_samp(26)  ), .I1 (px3202), .I2 (
         px3187), .I3 (px2953), .I4 (px2828), .I5 (px2641)) ;
         defparam ix19892z39819.INIT = 64'h9669699669969669;
    LUT6 ix19890z28344 (.O (px2642), .I0 (\p_key_samp(62)  ), .I1 (px3207), .I2 (
         px3206), .I3 (px3006), .I4 (px2857), .I5 (px2673)) ;
         defparam ix19890z28344.INIT = 64'h6996966996696996;
    LUT6 ix19889z39819 (.O (px2643), .I0 (\p_key_samp(29)  ), .I1 (px3217), .I2 (
         px3216), .I3 (px3010), .I4 (px2855), .I5 (px2671)) ;
         defparam ix19889z39819.INIT = 64'h9669699669969669;
    LUT6 ix19888z28344 (.O (px2644), .I0 (\p_key_samp(53)  ), .I1 (px3192), .I2 (
         px3191), .I3 (px3035), .I4 (px2836), .I5 (px2645)) ;
         defparam ix19888z28344.INIT = 64'h6996966996696996;
    LUT6 ix19886z39819 (.O (px2646), .I0 (\p_key_samp(39)  ), .I1 (px3198), .I2 (
         px3197), .I3 (px3054), .I4 (px2832), .I5 (px2647)) ;
         defparam ix19886z39819.INIT = 64'h9669699669969669;
    LUT6 ix18891z39819 (.O (px2654), .I0 (\p_key_samp(2)  ), .I1 (px3230), .I2 (
         px3229), .I3 (px2970), .I4 (px2818), .I5 (px2655)) ;
         defparam ix18891z39819.INIT = 64'h9669699669969669;
    LUT6 ix18889z28344 (.O (px2656), .I0 (\p_key_samp(52)  ), .I1 (px3227), .I2 (
         px3226), .I3 (px2967), .I4 (px2822), .I5 (px2657)) ;
         defparam ix18889z28344.INIT = 64'h6996966996696996;
    LUT6 ix18887z39819 (.O (px2658), .I0 (\p_key_samp(3)  ), .I1 (px3236), .I2 (
         px3235), .I3 (px2982), .I4 (px2824), .I5 (px2659)) ;
         defparam ix18887z39819.INIT = 64'h9669699669969669;
    LUT6 ix17894z28344 (.O (px2664), .I0 (\p_key_samp(9)  ), .I1 (px3233), .I2 (
         px3232), .I3 (px2973), .I4 (px2820), .I5 (px2665)) ;
         defparam ix17894z28344.INIT = 64'h6996966996696996;
    LUT6 ix17890z39819 (.O (px2668), .I0 (\p_key_samp(4)  ), .I1 (px3311), .I2 (
         px3296), .I3 (px3060), .I4 (px2893), .I5 (px2720)) ;
         defparam ix17890z39819.INIT = 64'h9669699669969669;
    LUT6 ix17889z39819 (.O (px2669), .I0 (\p_key_samp(28)  ), .I1 (px3294), .I2 (
         px3283), .I3 (px3077), .I4 (px2871), .I5 (px2710)) ;
         defparam ix17889z39819.INIT = 64'h9669699669969669;
    LUT6 ix16901z39819 (.O (px2670), .I0 (\p_key_samp(13)  ), .I1 (px3217), .I2 (
         px3216), .I3 (px3010), .I4 (px2855), .I5 (px2671)) ;
         defparam ix16901z39819.INIT = 64'h9669699669969669;
    LUT6 ix16899z28344 (.O (px2672), .I0 (\p_key_samp(55)  ), .I1 (px3207), .I2 (
         px3206), .I3 (px3006), .I4 (px2857), .I5 (px2673)) ;
         defparam ix16899z28344.INIT = 64'h6996966996696996;
    LUT6 ix16893z39819 (.O (px2678), .I0 (\p_key_samp(44)  ), .I1 (px3280), .I2 (
         px3245), .I3 (px2985), .I4 (px2790), .I5 (px2679)) ;
         defparam ix16893z39819.INIT = 64'h9669699669969669;
    LUT6 ix15904z39819 (.O (px2680), .I0 (\p_key_samp(50)  ), .I1 (px3262), .I2 (
         px3261), .I3 (px2987), .I4 (px2795), .I5 (px2681)) ;
         defparam ix15904z39819.INIT = 64'h9669699669969669;
    LUT6 ix15902z39819 (.O (px2682), .I0 (\p_key_samp(44)  ), .I1 (px3349), .I2 (
         px3330), .I3 (px3136), .I4 (px2927), .I5 (px2766)) ;
         defparam ix15902z39819.INIT = 64'h9669699669969669;
    LUT6 ix15901z39819 (.O (px2683), .I0 (\p_key_samp(1)  ), .I1 (px3328), .I2 (
         px3313), .I3 (px3090), .I4 (px2881), .I5 (px2732)) ;
         defparam ix15901z39819.INIT = 64'h9669699669969669;
    LUT6 ix14903z28344 (.O (px2694), .I0 (\p_key_samp(18)  ), .I1 (px3279), .I2 (
         px3278), .I3 (px2997), .I4 (px2798), .I5 (px2695)) ;
         defparam ix14903z28344.INIT = 64'h6996966996696996;
    LUT6 ix14899z28344 (.O (px2698), .I0 (\p_key_samp(6)  ), .I1 (px3308), .I2 (
         px3307), .I3 (px3073), .I4 (px2895), .I5 (px2728)) ;
         defparam ix14899z28344.INIT = 64'h6996966996696996;
    LUT6 ix12909z28344 (.O (px2702), .I0 (\p_key_samp(28)  ), .I1 (px3354), .I2 (
         px3353), .I3 (px3109), .I4 (px2907), .I5 (px2746)) ;
         defparam ix12909z28344.INIT = 64'h6996966996696996;
    LUT6 ix12908z28344 (.O (px2703), .I0 (\p_key_samp(61)  ), .I1 (px3374), .I2 (
         px3373), .I3 (px3112), .I4 (px2909), .I5 (px2752)) ;
         defparam ix12908z28344.INIT = 64'h6996966996696996;
    LUT6 ix12905z39819 (.O (px2706), .I0 (\p_key_samp(51)  ), .I1 (px3222), .I2 (
         px3221), .I3 (px3057), .I4 (px2868), .I5 (px2707)) ;
         defparam ix12905z39819.INIT = 64'h9669699669969669;
    LUT6 ix12902z39819 (.O (px2709), .I0 (\p_key_samp(12)  ), .I1 (px3294), .I2 (
         px3283), .I3 (px3077), .I4 (px2871), .I5 (px2710)) ;
         defparam ix12902z39819.INIT = 64'h9669699669969669;
    LUT6 ix11913z39819 (.O (px2711), .I0 (\p_key_samp(50)  ), .I1 (px3342), .I2 (
         px3341), .I3 (px3138), .I4 (px2929), .I5 (px2772)) ;
         defparam ix11913z39819.INIT = 64'h9669699669969669;
    LUT6 ix11912z39819 (.O (px2712), .I0 (\p_key_samp(36)  ), .I1 (px3444), .I2 (
         px3425), .I3 (px3170), .I4 (px3017), .I5 (px2802)) ;
         defparam ix11912z39819.INIT = 64'h9669699669969669;
    LUT6 ix11905z39819 (.O (px2719), .I0 (\p_key_samp(15)  ), .I1 (px3311), .I2 (
         px3296), .I3 (px3060), .I4 (px2893), .I5 (px2720)) ;
         defparam ix11905z39819.INIT = 64'h9669699669969669;
    LUT6 ix10914z28344 (.O (px2723), .I0 (\p_key_samp(2)  ), .I1 (px3333), .I2 (
         px3332), .I3 (px3154), .I4 (px2943), .I5 (px2770)) ;
         defparam ix10914z28344.INIT = 64'h6996966996696996;
    LUT6 ix10908z39819 (.O (px2729), .I0 (\p_key_samp(52)  ), .I1 (px3305), .I2 (
         px3304), .I3 (px3068), .I4 (px2899), .I5 (px2730)) ;
         defparam ix10908z39819.INIT = 64'h9669699669969669;
    LUT6 ix9919z39819 (.O (px2731), .I0 (\p_key_samp(46)  ), .I1 (px3328), .I2 (
         px3313), .I3 (px3090), .I4 (px2881), .I5 (px2732)) ;
         defparam ix9919z39819.INIT = 64'h9669699669969669;
    LUT6 ix9917z28344 (.O (px2733), .I0 (\p_key_samp(22)  ), .I1 (px3322), .I2 (
         px3321), .I3 (px3095), .I4 (px2885), .I5 (px2734)) ;
         defparam ix9917z28344.INIT = 64'h6996966996696996;
    LUT6 ix8922z28344 (.O (px2741), .I0 (\p_key_samp(15)  ), .I1 (px3316), .I2 (
         px3315), .I3 (px3092), .I4 (px2891), .I5 (px2742)) ;
         defparam ix8922z28344.INIT = 64'h6996966996696996;
    LUT6 ix7925z28344 (.O (px2751), .I0 (\p_key_samp(12)  ), .I1 (px3374), .I2 (
         px3373), .I3 (px3112), .I4 (px2909), .I5 (px2752)) ;
         defparam ix7925z28344.INIT = 64'h6996966996696996;
    LUT6 ix6929z39819 (.O (px2760), .I0 (\p_key_samp(52)  ), .I1 (px3411), .I2 (
         px3410), .I3 (px3261), .I4 (px2987), .I5 (px2795)) ;
         defparam ix6929z39819.INIT = 64'h9669699669969669;
    LUT6 ix6926z28344 (.O (px2763), .I0 (\p_key_samp(42)  ), .I1 (px3452), .I2 (
         px3451), .I3 (px3235), .I4 (px2982), .I5 (px2824)) ;
         defparam ix6926z28344.INIT = 64'h6996966996696996;
    LUT6 ix6925z28344 (.O (px2764), .I0 (\p_key_samp(39)  ), .I1 (px3723), .I2 (
         px3504), .I3 (px3281), .I4 (px3058), .I5 (px2869)) ;
         defparam ix6925z28344.INIT = 64'h6996966996696996;
    LUT6 ix6924z39819 (.O (px2765), .I0 (\p_key_samp(22)  ), .I1 (px3349), .I2 (
         px3330), .I3 (px3136), .I4 (px2927), .I5 (px2766)) ;
         defparam ix6924z39819.INIT = 64'h9669699669969669;
    LUT6 ix5929z39819 (.O (px2773), .I0 (\p_key_samp(3)  ), .I1 (px3434), .I2 (
         px3433), .I3 (px3183), .I4 (px3041), .I5 (px2811)) ;
         defparam ix5929z39819.INIT = 64'h9669699669969669;
    LUT6 ix5925z39819 (.O (px2777), .I0 (\p_key_samp(26)  ), .I1 (px3455), .I2 (
         px3454), .I3 (px3226), .I4 (px2967), .I5 (px2822)) ;
         defparam ix5925z39819.INIT = 64'h9669699669969669;
    LUT6 ix4935z28344 (.O (px2780), .I0 (\p_key_samp(41)  ), .I1 (px3440), .I2 (
         px3439), .I3 (px3172), .I4 (px3022), .I5 (px2807)) ;
         defparam ix4935z28344.INIT = 64'h6996966996696996;
    LUT6 ix3935z28344 (.O (px2793), .I0 (\p_key_samp(43)  ), .I1 (px3551), .I2 (
         px3536), .I3 (px3330), .I4 (px3136), .I5 (px2927)) ;
         defparam ix3935z28344.INIT = 64'h6996966996696996;
    LUT6 ix3934z39819 (.O (px2794), .I0 (\p_key_samp(18)  ), .I1 (px3411), .I2 (
         px3410), .I3 (px3261), .I4 (px2987), .I5 (px2795)) ;
         defparam ix3934z39819.INIT = 64'h9669699669969669;
    LUT6 ix3932z39819 (.O (px2796), .I0 (\p_key_samp(36)  ), .I1 (px3521), .I2 (
         px3506), .I3 (px3313), .I4 (px3090), .I5 (px2881)) ;
         defparam ix3932z39819.INIT = 64'h9669699669969669;
    LUT6 ix3931z28344 (.O (px2797), .I0 (\p_key_samp(49)  ), .I1 (px3422), .I2 (
         px3421), .I3 (px3278), .I4 (px2997), .I5 (px2798)) ;
         defparam ix3931z28344.INIT = 64'h6996966996696996;
    LUT6 ix1941z39819 (.O (px2801), .I0 (\p_key_samp(42)  ), .I1 (px3444), .I2 (
         px3425), .I3 (px3170), .I4 (px3017), .I5 (px2802)) ;
         defparam ix1941z39819.INIT = 64'h9669699669969669;
    LUT6 ix1939z28344 (.O (px2803), .I0 (\p_key_samp(6)  ), .I1 (px3443), .I2 (
         px3442), .I3 (px3191), .I4 (px3035), .I5 (px2836)) ;
         defparam ix1939z28344.INIT = 64'h6996966996696996;
    LUT6 ix945z39819 (.O (px2810), .I0 (\p_key_samp(53)  ), .I1 (px3434), .I2 (
         px3433), .I3 (px3183), .I4 (px3041), .I5 (px2811)) ;
         defparam ix945z39819.INIT = 64'h9669699669969669;
    LUT6 ix943z28344 (.O (px2812), .I0 (\p_key_samp(28)  ), .I1 (px3437), .I2 (
         px3436), .I3 (px3197), .I4 (px3054), .I5 (px2832)) ;
         defparam ix943z28344.INIT = 64'h6996966996696996;
    LUT6 ix65483z39819 (.O (px2821), .I0 (\p_key_samp(51)  ), .I1 (px3455), .I2 (
         px3454), .I3 (px3226), .I4 (px2967), .I5 (px2822)) ;
         defparam ix65483z39819.INIT = 64'h9669699669969669;
    LUT6 ix65481z28344 (.O (px2823), .I0 (\p_key_samp(34)  ), .I1 (px3452), .I2 (
         px3451), .I3 (px3235), .I4 (px2982), .I5 (px2824)) ;
         defparam ix65481z28344.INIT = 64'h6996966996696996;
    LUT6 ix65477z39819 (.O (px2827), .I0 (\p_key_samp(57)  ), .I1 (px3403), .I2 (
         px3392), .I3 (px3187), .I4 (px2953), .I5 (px2828)) ;
         defparam ix65477z39819.INIT = 64'h9669699669969669;
    LUT6 ix64482z28344 (.O (px2835), .I0 (\p_key_samp(21)  ), .I1 (px3443), .I2 (
         px3442), .I3 (px3191), .I4 (px3035), .I5 (px2836)) ;
         defparam ix64482z28344.INIT = 64'h6996966996696996;
    LUT6 ix63489z28344 (.O (px2841), .I0 (\p_key_samp(37)  ), .I1 (px3611), .I2 (
         px3582), .I3 (px3296), .I4 (px3060), .I5 (px2893)) ;
         defparam ix63489z28344.INIT = 64'h6996966996696996;
    LUT6 ix63486z28344 (.O (px2844), .I0 (\p_key_samp(14)  ), .I1 (px3886), .I2 (
         px3724), .I3 (px3504), .I4 (px3281), .I5 (px3058)) ;
         defparam ix63486z28344.INIT = 64'h6996966996696996;
    LUT6 ix63485z39819 (.O (px2845), .I0 (\p_key_samp(46)  ), .I1 (px3576), .I2 (
         px3565), .I3 (px3359), .I4 (px3119), .I5 (px2914)) ;
         defparam ix63485z39819.INIT = 64'h9669699669969669;
    LUT6 ix63484z28344 (.O (px2846), .I0 (\p_key_samp(5)  ), .I1 (px3512), .I2 (
         px3511), .I3 (px3321), .I4 (px3095), .I5 (px2885)) ;
         defparam ix63484z28344.INIT = 64'h6996966996696996;
    LUT6 ix63483z28344 (.O (px2847), .I0 (\p_key_samp(20)  ), .I1 (px3515), .I2 (
         px3514), .I3 (px3315), .I4 (px3092), .I5 (px2891)) ;
         defparam ix63483z28344.INIT = 64'h6996966996696996;
    LUT6 ix62485z39819 (.O (px2858), .I0 (\p_key_samp(29)  ), .I1 (px3563), .I2 (
         px3562), .I3 (px3373), .I4 (px3112), .I5 (px2909)) ;
         defparam ix62485z39819.INIT = 64'h9669699669969669;
    LUT6 ix62484z28344 (.O (px2859), .I0 (\p_key_samp(61)  ), .I1 (px3560), .I2 (
         px3559), .I3 (px3353), .I4 (px3109), .I5 (px2907)) ;
         defparam ix62484z28344.INIT = 64'h6996966996696996;
    LUT6 ix61496z28344 (.O (px2860), .I0 (\p_key_samp(63)  ), .I1 (px3588), .I2 (
         px3587), .I3 (px3304), .I4 (px3068), .I5 (px2899)) ;
         defparam ix61496z28344.INIT = 64'h6996966996696996;
    LUT6 ix61491z28344 (.O (px2865), .I0 (\p_key_samp(39)  ), .I1 (px3607), .I2 (
         px3596), .I3 (px3307), .I4 (px3073), .I5 (px2895)) ;
         defparam ix61491z28344.INIT = 64'h6996966996696996;
    LUT6 ix61490z39819 (.O (px2866), .I0 (\p_key_samp(61)  ), .I1 (px3534), .I2 (
         px3523), .I3 (px3283), .I4 (px3077), .I5 (px2871)) ;
         defparam ix61490z39819.INIT = 64'h9669699669969669;
    LUT6 ix61489z39819 (.O (px2867), .I0 (\p_key_samp(19)  ), .I1 (px3406), .I2 (
         px3405), .I3 (px3221), .I4 (px3057), .I5 (px2868)) ;
         defparam ix61489z39819.INIT = 64'h9669699669969669;
    LUT6 ix60499z39819 (.O (px2870), .I0 (\p_key_samp(45)  ), .I1 (px3534), .I2 (
         px3523), .I3 (px3283), .I4 (px3077), .I5 (px2871)) ;
         defparam ix60499z39819.INIT = 64'h9669699669969669;
    LUT6 ix60497z28344 (.O (px2872), .I0 (\p_key_samp(18)  ), .I1 (px3544), .I2 (
         px3543), .I3 (px3341), .I4 (px3138), .I5 (px2929)) ;
         defparam ix60497z28344.INIT = 64'h6996966996696996;
    LUT6 ix60492z28344 (.O (px2877), .I0 (\p_key_samp(35)  ), .I1 (px3630), .I2 (
         px3615), .I3 (px3425), .I4 (px3170), .I5 (px3017)) ;
         defparam ix60492z28344.INIT = 64'h6996966996696996;
    LUT6 ix60491z28344 (.O (px2878), .I0 (\p_key_samp(17)  ), .I1 (px3667), .I2 (
         px3652), .I3 (px3408), .I4 (px3245), .I5 (px2985)) ;
         defparam ix60491z28344.INIT = 64'h6996966996696996;
    LUT6 ix60490z39819 (.O (px2879), .I0 (\p_key_samp(59)  ), .I1 (px3547), .I2 (
         px3546), .I3 (px3338), .I4 (px3160), .I5 (px2945)) ;
         defparam ix60490z39819.INIT = 64'h9669699669969669;
    LUT6 ix59498z28344 (.O (px2884), .I0 (\p_key_samp(55)  ), .I1 (px3512), .I2 (
         px3511), .I3 (px3321), .I4 (px3095), .I5 (px2885)) ;
         defparam ix59498z28344.INIT = 64'h6996966996696996;
    LUT6 ix59496z28344 (.O (px2886), .I0 (\p_key_samp(31)  ), .I1 (px3647), .I2 (
         px3632), .I3 (px3392), .I4 (px3187), .I5 (px2953)) ;
         defparam ix59496z28344.INIT = 64'h6996966996696996;
    LUT6 ix59495z39819 (.O (px2887), .I0 (\p_key_samp(37)  ), .I1 (px3650), .I2 (
         px3649), .I3 (px3405), .I4 (px3221), .I5 (px3057)) ;
         defparam ix59495z39819.INIT = 64'h9669699669969669;
    LUT6 ix58505z28344 (.O (px2890), .I0 (\p_key_samp(12)  ), .I1 (px3515), .I2 (
         px3514), .I3 (px3315), .I4 (px3092), .I5 (px2891)) ;
         defparam ix58505z28344.INIT = 64'h6996966996696996;
    LUT6 ix58503z28344 (.O (px2892), .I0 (\p_key_samp(12)  ), .I1 (px3611), .I2 (
         px3582), .I3 (px3296), .I4 (px3060), .I5 (px2893)) ;
         defparam ix58503z28344.INIT = 64'h6996966996696996;
    LUT6 ix58501z28344 (.O (px2894), .I0 (\p_key_samp(27)  ), .I1 (px3607), .I2 (
         px3596), .I3 (px3307), .I4 (px3073), .I5 (px2895)) ;
         defparam ix58501z28344.INIT = 64'h6996966996696996;
    LUT6 ix58499z28344 (.O (px2896), .I0 (\p_key_samp(2)  ), .I1 (px3591), .I2 (
         px3590), .I3 (px3335), .I4 (px3151), .I5 (px2941)) ;
         defparam ix58499z28344.INIT = 64'h6996966996696996;
    LUT6 ix58498z28344 (.O (px2897), .I0 (\p_key_samp(33)  ), .I1 (px3585), .I2 (
         px3584), .I3 (px3332), .I4 (px3154), .I5 (px2943)) ;
         defparam ix58498z28344.INIT = 64'h6996966996696996;
    LUT6 ix58497z28344 (.O (px2898), .I0 (\p_key_samp(51)  ), .I1 (px3588), .I2 (
         px3587), .I3 (px3304), .I4 (px3068), .I5 (px2899)) ;
         defparam ix58497z28344.INIT = 64'h6996966996696996;
    LUT6 ix56503z28344 (.O (px2906), .I0 (\p_key_samp(21)  ), .I1 (px3560), .I2 (
         px3559), .I3 (px3353), .I4 (px3109), .I5 (px2907)) ;
         defparam ix56503z28344.INIT = 64'h6996966996696996;
    LUT6 ix56501z39819 (.O (px2908), .I0 (\p_key_samp(45)  ), .I1 (px3563), .I2 (
         px3562), .I3 (px3373), .I4 (px3112), .I5 (px2909)) ;
         defparam ix56501z39819.INIT = 64'h9669699669969669;
    LUT6 ix55510z28344 (.O (px2912), .I0 (\p_key_samp(7)  ), .I1 (px3886), .I2 (
         px3724), .I3 (px3504), .I4 (px3281), .I5 (px3058)) ;
         defparam ix55510z28344.INIT = 64'h6996966996696996;
    LUT6 ix55509z39819 (.O (px2913), .I0 (\p_key_samp(30)  ), .I1 (px3576), .I2 (
         px3565), .I3 (px3359), .I4 (px3119), .I5 (px2914)) ;
         defparam ix55509z39819.INIT = 64'h9669699669969669;
    LUT6 ix54514z28344 (.O (px2921), .I0 (\p_key_samp(42)  ), .I1 (px3666), .I2 (
         px3665), .I3 (px3421), .I4 (px3278), .I5 (px2997)) ;
         defparam ix54514z28344.INIT = 64'h6996966996696996;
    LUT6 ix54511z28344 (.O (px2924), .I0 (\p_key_samp(51)  ), .I1 (px3658), .I2 (
         px3657), .I3 (px3410), .I4 (px3261), .I5 (px2987)) ;
         defparam ix54511z28344.INIT = 64'h6996966996696996;
    LUT6 ix54510z28344 (.O (px2925), .I0 (\p_key_samp(10)  ), .I1 (px3703), .I2 (
         px3702), .I3 (px3451), .I4 (px3235), .I5 (px2982)) ;
         defparam ix54510z28344.INIT = 64'h6996966996696996;
    LUT6 ix54509z28344 (.O (px2926), .I0 (\p_key_samp(55)  ), .I1 (px3551), .I2 (
         px3536), .I3 (px3330), .I4 (px3136), .I5 (px2927)) ;
         defparam ix54509z28344.INIT = 64'h6996966996696996;
    LUT6 ix54507z28344 (.O (px2928), .I0 (\p_key_samp(26)  ), .I1 (px3544), .I2 (
         px3543), .I3 (px3341), .I4 (px3138), .I5 (px2929)) ;
         defparam ix54507z28344.INIT = 64'h6996966996696996;
    LUT6 ix53515z39819 (.O (px2933), .I0 (\p_key_samp(9)  ), .I1 (px3624), .I2 (
         px3623), .I3 (px3439), .I4 (px3172), .I5 (px3022)) ;
         defparam ix53515z39819.INIT = 64'h9669699669969669;
    LUT6 ix53514z28344 (.O (px2934), .I0 (\p_key_samp(34)  ), .I1 (px3627), .I2 (
         px3626), .I3 (px3433), .I4 (px3183), .I5 (px3041)) ;
         defparam ix53514z28344.INIT = 64'h6996966996696996;
    LUT6 ix53513z28344 (.O (px2935), .I0 (\p_key_samp(57)  ), .I1 (px3717), .I2 (
         px3716), .I3 (px3454), .I4 (px3226), .I5 (px2967)) ;
         defparam ix53513z28344.INIT = 64'h6996966996696996;
    LUT6 ix53509z39819 (.O (px2939), .I0 (\p_key_samp(58)  ), .I1 (px3689), .I2 (
         px3688), .I3 (px3448), .I4 (px3229), .I5 (px2970)) ;
         defparam ix53509z39819.INIT = 64'h9669699669969669;
    LUT6 ix52521z28344 (.O (px2940), .I0 (\p_key_samp(36)  ), .I1 (px3591), .I2 (
         px3590), .I3 (px3335), .I4 (px3151), .I5 (px2941)) ;
         defparam ix52521z28344.INIT = 64'h6996966996696996;
    LUT6 ix52519z28344 (.O (px2942), .I0 (\p_key_samp(58)  ), .I1 (px3585), .I2 (
         px3584), .I3 (px3332), .I4 (px3154), .I5 (px2943)) ;
         defparam ix52519z28344.INIT = 64'h6996966996696996;
    LUT6 ix52517z39819 (.O (px2944), .I0 (\p_key_samp(49)  ), .I1 (px3547), .I2 (
         px3546), .I3 (px3338), .I4 (px3160), .I5 (px2945)) ;
         defparam ix52517z39819.INIT = 64'h9669699669969669;
    LUT6 ix51522z28344 (.O (px2952), .I0 (\p_key_samp(25)  ), .I1 (px3647), .I2 (
         px3632), .I3 (px3392), .I4 (px3187), .I5 (px2953)) ;
         defparam ix51522z28344.INIT = 64'h6996966996696996;
    LUT6 ix51515z28344 (.O (px2959), .I0 (\p_key_samp(63)  ), .I1 (px3675), .I2 (
         px3674), .I3 (px3483), .I4 (px3206), .I5 (px3006)) ;
         defparam ix51515z28344.INIT = 64'h6996966996696996;
    LUT6 ix50524z28344 (.O (px2963), .I0 (\p_key_samp(54)  ), .I1 (px3639), .I2 (
         px3638), .I3 (px3442), .I4 (px3191), .I5 (px3035)) ;
         defparam ix50524z28344.INIT = 64'h6996966996696996;
    LUT6 ix50521z28344 (.O (px2966), .I0 (\p_key_samp(19)  ), .I1 (px3717), .I2 (
         px3716), .I3 (px3454), .I4 (px3226), .I5 (px2967)) ;
         defparam ix50521z28344.INIT = 64'h6996966996696996;
    LUT6 ix50518z39819 (.O (px2969), .I0 (\p_key_samp(1)  ), .I1 (px3689), .I2 (
         px3688), .I3 (px3448), .I4 (px3229), .I5 (px2970)) ;
         defparam ix50518z39819.INIT = 64'h9669699669969669;
    LUT6 ix49528z39819 (.O (px2972), .I0 (\p_key_samp(43)  ), .I1 (px3714), .I2 (
         px3705), .I3 (px3460), .I4 (px3232), .I5 (px2973)) ;
         defparam ix49528z39819.INIT = 64'h9669699669969669;
    LUT6 ix48532z28344 (.O (px2981), .I0 (\p_key_samp(2)  ), .I1 (px3703), .I2 (
         px3702), .I3 (px3451), .I4 (px3235), .I5 (px2982)) ;
         defparam ix48532z28344.INIT = 64'h6996966996696996;
    LUT6 ix48529z28344 (.O (px2984), .I0 (\p_key_samp(11)  ), .I1 (px3667), .I2 (
         px3652), .I3 (px3408), .I4 (px3245), .I5 (px2985)) ;
         defparam ix48529z28344.INIT = 64'h6996966996696996;
    LUT6 ix48527z28344 (.O (px2986), .I0 (\p_key_samp(49)  ), .I1 (px3658), .I2 (
         px3657), .I3 (px3410), .I4 (px3261), .I5 (px2987)) ;
         defparam ix48527z28344.INIT = 64'h6996966996696996;
    LUT6 ix47530z28344 (.O (px2996), .I0 (\p_key_samp(17)  ), .I1 (px3666), .I2 (
         px3665), .I3 (px3421), .I4 (px3278), .I5 (px2997)) ;
         defparam ix47530z28344.INIT = 64'h6996966996696996;
    LUT6 ix47527z39819 (.O (px2999), .I0 (\p_key_samp(35)  ), .I1 (px3750), .I2 (
         px3739), .I3 (px3506), .I4 (px3313), .I5 (px3090)) ;
         defparam ix47527z39819.INIT = 64'h9669699669969669;
    LUT6 ix32964z28344 (.O (px3005), .I0 (\p_key_samp(20)  ), .I1 (px3675), .I2 (
         px3674), .I3 (px3483), .I4 (px3206), .I5 (px3006)) ;
         defparam ix32964z28344.INIT = 64'h6996966996696996;
    LUT6 ix32967z28344 (.O (px3008), .I0 (\p_key_samp(5)  ), .I1 (px3737), .I2 (
         px3726), .I3 (px3582), .I4 (px3296), .I5 (px3060)) ;
         defparam ix32967z28344.INIT = 64'h6996966996696996;
    LUT6 ix33961z39819 (.O (px3015), .I0 (\p_key_samp(29)  ), .I1 (px3761), .I2 (
         px3752), .I3 (px3523), .I4 (px3283), .I5 (px3077)) ;
         defparam ix33961z39819.INIT = 64'h9669699669969669;
    LUT6 ix33962z28344 (.O (px3016), .I0 (\p_key_samp(10)  ), .I1 (px3630), .I2 (
         px3615), .I3 (px3425), .I4 (px3170), .I5 (px3017)) ;
         defparam ix33962z28344.INIT = 64'h6996966996696996;
    LUT6 ix34954z39819 (.O (px3021), .I0 (\p_key_samp(15)  ), .I1 (px3624), .I2 (
         px3623), .I3 (px3439), .I4 (px3172), .I5 (px3022)) ;
         defparam ix34954z39819.INIT = 64'h9669699669969669;
    LUT6 ix35954z28344 (.O (px3034), .I0 (\p_key_samp(39)  ), .I1 (px3639), .I2 (
         px3638), .I3 (px3442), .I4 (px3191), .I5 (px3035)) ;
         defparam ix35954z28344.INIT = 64'h6996966996696996;
    LUT6 ix36947z28344 (.O (px3040), .I0 (\p_key_samp(21)  ), .I1 (px3627), .I2 (
         px3626), .I3 (px3433), .I4 (px3183), .I5 (px3041)) ;
         defparam ix36947z28344.INIT = 64'h6996966996696996;
    LUT6 ix37947z28344 (.O (px3053), .I0 (\p_key_samp(61)  ), .I1 (px3636), .I2 (
         px3635), .I3 (px3436), .I4 (px3197), .I5 (px3054)) ;
         defparam ix37947z28344.INIT = 64'h6996966996696996;
    LUT6 ix37950z39819 (.O (px3056), .I0 (\p_key_samp(50)  ), .I1 (px3650), .I2 (
         px3649), .I3 (px3405), .I4 (px3221), .I5 (px3057)) ;
         defparam ix37950z39819.INIT = 64'h9669699669969669;
    LUT6 ix37953z28344 (.O (px3059), .I0 (\p_key_samp(45)  ), .I1 (px3737), .I2 (
         px3726), .I3 (px3582), .I4 (px3296), .I5 (px3060)) ;
         defparam ix37953z28344.INIT = 64'h6996966996696996;
    LUT6 ix39944z39819 (.O (px3076), .I0 (\p_key_samp(13)  ), .I1 (px3761), .I2 (
         px3752), .I3 (px3523), .I4 (px3283), .I5 (px3077)) ;
         defparam ix39944z39819.INIT = 64'h9669699669969669;
    LUT6 ix40944z39819 (.O (px3089), .I0 (\p_key_samp(47)  ), .I1 (px3750), .I2 (
         px3739), .I3 (px3506), .I4 (px3313), .I5 (px3090)) ;
         defparam ix40944z39819.INIT = 64'h9669699669969669;
    LUT3 ix42217z1464 (.O (px3697), .I0 (\p_plaintext(39)  ), .I1 (
         \p_key_samp(6)  ), .I2 (px3781)) ;
         defparam ix42217z1464.INIT = 8'h96;
    LUT3 ix48198z1464 (.O (px3744), .I0 (\p_plaintext(37)  ), .I1 (
         \p_key_samp(22)  ), .I2 (px3745)) ;
         defparam ix48198z1464.INIT = 8'h96;
    LUT2 ix62154z1320 (.O (px3870), .I0 (\p_plaintext(63)  ), .I1 (
         \p_key_samp(61)  )) ;
         defparam ix62154z1320.INIT = 4'h6;
    LUT2 ix62156z1320 (.O (px3872), .I0 (\p_plaintext(37)  ), .I1 (
         \p_key_samp(6)  )) ;
         defparam ix62156z1320.INIT = 4'h6;
    LUT2 ix2605z1320 (.O (px3923), .I0 (\p_plaintext(5)  ), .I1 (
         \p_key_samp(22)  )) ;
         defparam ix2605z1320.INIT = 4'h6;
endmodule


module input_register_0 ( px3886, px3870, px3872, px3923, px3761, px3750, px3737, 
                          px3717, px3703, px3689, px3675, px3667, px3666, px3658, 
                          px3650, px3647, px3639, px3630, px3627, px3697, px3624, 
                          px3611, px3607, px3744, px3591, px3588, px3585, px3576, 
                          px3563, px3560, px3551, px3547, px3544, px3534, px3515, 
                          px3512, px3455, px3452, px3444, px3443, px3434, px3411, 
                          px3374, px3739, px3649, px3632, px3523, px3752, px3652, 
                          px3546, px3425, px3615, px3543, px3582, px3726, px3584, 
                          px3590, px3433, px3626, px3596, px3587, px3559, px3781, 
                          px3373, px3562, px3442, px3638, px3623, px3511, px3514, 
                          px3745, px3724, px3565, px3674, px3665, px3536, px3410, 
                          px3657, px3451, px3702, px3688, px3454, px3716, px3635, 
                          px3636, px3705, px3714, px2959, px2963, px2986, px2996, 
                          px2999, px3506, px3521, px3089, px3059, px3076, px2921, 
                          px2925, px2924, px2933, px2934, px2935, px2939, px3005, 
                          px3008, px3015, \p_key_samp(15)  , px2966, px2969, 
                          px2972, px2981, px3021, px3034, px3040, px3053, px3436, 
                          px3437, px3483, px2928, px2944, px2942, px2940, 
                          \p_key_samp(44)  , px2952, px2984, px3016, px3056, 
                          px3439, px3440, px2865, px2859, px2858, px2860, px2844, 
                          px2845, px2846, px2847, \p_key_samp(50)  , px2872, 
                          px2877, px2878, px2879, px3448, px2912, px2908, px2906, 
                          px2913, px3341, px3342, px3332, px3333, px2894, px2896, 
                          px2897, px2898, px2884, px2886, px2887, px2890, px3421, 
                          px3422, px3460, px3353, px3354, px3405, px3406, 
                          \p_key_samp(4)  , px3392, px3403, px2793, px2794, 
                          px2796, px2797, \p_key_samp(45)  , px3307, px3308, 
                          px3335, px2835, px3408, px3338, px2763, px2760, px2892, 
                          px2870, px2926, px2773, px2777, px2780, px3304, px3305, 
                          px2841, px2866, px2821, px2823, px3359, 
                          \p_key_samp(13)  , px3504, px3723, px3315, px3316, 
                          px3321, px3322, px2803, px2810, px2812, 
                          \p_key_samp(6)  , px2801, px2867, px2827, px2698, 
                          px2702, px2703, \p_key_samp(61)  , px2733, px2741, 
                          px2723, px2729, px2711, px2712, px2764, px2751, 
                          \p_key_samp(10)  , \p_key_samp(46)  , px2680, px2682, 
                          px2683, px2694, \p_key_samp(21)  , \p_key_samp(12)  , 
                          \p_key_samp(5)  , \p_key_samp(7)  , px2765, px2719, 
                          px2709, px2731, \p_key_samp(49)  , px2642, px2643, 
                          px2644, px2646, px2618, px2621, px2622, px2623, 
                          \p_key_samp(39)  , \p_key_samp(47)  , \p_key_samp(28)  , 
                          px2654, px2656, px2658, px2664, \p_key_samp(23)  , 
                          px2630, px2634, px2637, px2638, \p_key_samp(22)  , 
                          \p_key_samp(54)  , \p_key_samp(37)  , px2668, px2670, 
                          px2669, px2672, px2605, px2606, px2607, px2608, px3007, 
                          \p_key_samp(14)  , \p_key_samp(63)  , \p_key_samp(30)  , 
                          \p_key_samp(53)  , \p_key_samp(31)  , px2514, px2507, 
                          \p_key_samp(29)  , \p_key_samp(20)  , px3036, 
                          \p_key_samp(62)  , \p_key_samp(38)  , \p_key_samp(55)  , 
                          px2497, \p_key_samp(19)  , \p_key_samp(52)  , px3052, 
                          \p_key_samp(59)  , \p_key_samp(34)  , \p_key_samp(2)  , 
                          \p_key_samp(17)  , \p_key_samp(26)  , px2585, px2591, 
                          px2587, px2593, \p_key_samp(51)  , \p_key_samp(3)  , 
                          \p_key_samp(33)  , \p_key_samp(9)  , px2628, px2640, 
                          px2678, px2706, \p_key_samp(27)  , \p_key_samp(35)  , 
                          \p_key_samp(58)  , px2570, px2569, px2566, px2563, 
                          \p_key_samp(36)  , px2573, px2575, px2579, px2582, 
                          \p_key_samp(18)  , px2601, px2611, px2613, px2615, 
                          \p_key_samp(41)  , px2551, px2555, px2557, px2558, 
                          \p_key_samp(60)  , \p_key_samp(25)  , \p_key_samp(42)  , 
                          \p_key_samp(1)  , \p_key_samp(11)  , px2528, px2523, 
                          px2522, px2521, \p_key_samp(57)  , px2537, px2534, 
                          px2533, px2538, \p_key_samp(43)  , px2708, px2869, 
                          px3058, px3281, px3503, px2432, px2707, px2868, px3057, 
                          px3221, px3222, px2431, px2430, px2429, px2576, px2742, 
                          px2891, px3092, px3093, px2428, px2588, px2768, px2941, 
                          px3151, px3152, px2427, px2426, px2425, px2592, px2786, 
                          px2945, px3160, px3161, px2424, px2641, px2828, px2953, 
                          px3187, px3202, px2423, px2422, px2421, px2420, px2629, 
                          px2802, px3017, px3170, px3185, px2419, px2418, px2556, 
                          px2730, px2899, px3068, px3069, px2417, px2602, px2748, 
                          px2914, px3119, px3120, px2416, px2415, px2594, px2772, 
                          px2929, px3138, px3149, px2414, px2413, px2614, px2752, 
                          px2909, px3112, px3113, px2412, px2586, px2770, px2943, 
                          px3154, px3155, px2411, px2410, px2409, px2552, px2728, 
                          px2895, px3073, px3074, px2408, px2574, px2734, px2885, 
                          px3095, px3096, px2407, px2406, px2405, px2612, px2746, 
                          px2907, px3109, px3110, px2404, px2403, px2402, px2679, 
                          px2790, px2985, px3245, px3280, px2401, px2671, px2855, 
                          px3010, px3216, px3217, px2400, px2639, px2807, px3022, 
                          px3172, px3173, px2399, px2665, px2820, px2973, px3232, 
                          px3233, px2398, px2766, px2927, px3136, px3330, px3349, 
                          px2397, px2396, px2395, px2394, px2393, px2392, px2391, 
                          px2390, px2389, px2720, px2893, px3060, px3296, px3311, 
                          px2388, px2647, px2832, px3054, px3197, px3198, px2387, 
                          px2655, px2818, px2970, px3229, px3230, px2386, px2695, 
                          px2798, px2997, px3278, px3279, px2385, px2710, px2871, 
                          px3077, px3283, px3294, px2384, px2508, px2645, px2836, 
                          px3035, px3191, px3192, px2383, px2657, px2822, px2967, 
                          px3226, px3227, px2382, px2681, px2795, px2987, px3261, 
                          px3262, px2381, px2380, px2379, px2378, px2377, px2376, 
                          px2375, px2374, px2373, px2732, px2881, px3090, px3313, 
                          px3328, px2372, px2520, px2673, px2857, px3006, px3206, 
                          px3207, px2371, px2498, px2631, px2811, px3041, px3183, 
                          px3184, px2370, px2659, px2824, px2982, px3235, px3236, 
                          px2369, p_nbus_data_in_int, p_nbus_plaintext, 
                          \p_plaintext(37)  , \p_plaintext(39)  , p_reset_int, 
                          p_load_int, p_clk_int, \p_plaintext(63)   ) ;

    output px3886 ;
    input px3870 ;
    input px3872 ;
    input px3923 ;
    output px3761 ;
    output px3750 ;
    output px3737 ;
    output px3717 ;
    output px3703 ;
    output px3689 ;
    output px3675 ;
    output px3667 ;
    output px3666 ;
    output px3658 ;
    output px3650 ;
    output px3647 ;
    output px3639 ;
    output px3630 ;
    output px3627 ;
    input px3697 ;
    output px3624 ;
    output px3611 ;
    output px3607 ;
    input px3744 ;
    output px3591 ;
    output px3588 ;
    output px3585 ;
    output px3576 ;
    output px3563 ;
    output px3560 ;
    output px3551 ;
    output px3547 ;
    output px3544 ;
    output px3534 ;
    output px3515 ;
    output px3512 ;
    output px3455 ;
    output px3452 ;
    output px3444 ;
    output px3443 ;
    output px3434 ;
    output px3411 ;
    output px3374 ;
    output px3739 ;
    output px3649 ;
    output px3632 ;
    output px3523 ;
    output px3752 ;
    output px3652 ;
    output px3546 ;
    output px3425 ;
    output px3615 ;
    output px3543 ;
    output px3582 ;
    output px3726 ;
    output px3584 ;
    output px3590 ;
    output px3433 ;
    output px3626 ;
    output px3596 ;
    output px3587 ;
    output px3559 ;
    output px3781 ;
    output px3373 ;
    output px3562 ;
    output px3442 ;
    output px3638 ;
    output px3623 ;
    output px3511 ;
    output px3514 ;
    output px3745 ;
    output px3724 ;
    output px3565 ;
    output px3674 ;
    output px3665 ;
    output px3536 ;
    output px3410 ;
    output px3657 ;
    output px3451 ;
    output px3702 ;
    output px3688 ;
    output px3454 ;
    output px3716 ;
    output px3635 ;
    output px3636 ;
    output px3705 ;
    output px3714 ;
    input px2959 ;
    input px2963 ;
    input px2986 ;
    input px2996 ;
    input px2999 ;
    output px3506 ;
    output px3521 ;
    input px3089 ;
    input px3059 ;
    input px3076 ;
    input px2921 ;
    input px2925 ;
    input px2924 ;
    input px2933 ;
    input px2934 ;
    input px2935 ;
    input px2939 ;
    input px3005 ;
    input px3008 ;
    input px3015 ;
    input \p_key_samp(15)   ;
    input px2966 ;
    input px2969 ;
    input px2972 ;
    input px2981 ;
    input px3021 ;
    input px3034 ;
    input px3040 ;
    input px3053 ;
    output px3436 ;
    output px3437 ;
    output px3483 ;
    input px2928 ;
    input px2944 ;
    input px2942 ;
    input px2940 ;
    input \p_key_samp(44)   ;
    input px2952 ;
    input px2984 ;
    input px3016 ;
    input px3056 ;
    output px3439 ;
    output px3440 ;
    input px2865 ;
    input px2859 ;
    input px2858 ;
    input px2860 ;
    input px2844 ;
    input px2845 ;
    input px2846 ;
    input px2847 ;
    input \p_key_samp(50)   ;
    input px2872 ;
    input px2877 ;
    input px2878 ;
    input px2879 ;
    output px3448 ;
    input px2912 ;
    input px2908 ;
    input px2906 ;
    input px2913 ;
    output px3341 ;
    output px3342 ;
    output px3332 ;
    output px3333 ;
    input px2894 ;
    input px2896 ;
    input px2897 ;
    input px2898 ;
    input px2884 ;
    input px2886 ;
    input px2887 ;
    input px2890 ;
    output px3421 ;
    output px3422 ;
    output px3460 ;
    output px3353 ;
    output px3354 ;
    output px3405 ;
    output px3406 ;
    input \p_key_samp(4)   ;
    output px3392 ;
    output px3403 ;
    input px2793 ;
    input px2794 ;
    input px2796 ;
    input px2797 ;
    input \p_key_samp(45)   ;
    output px3307 ;
    output px3308 ;
    output px3335 ;
    input px2835 ;
    output px3408 ;
    output px3338 ;
    input px2763 ;
    input px2760 ;
    input px2892 ;
    input px2870 ;
    input px2926 ;
    input px2773 ;
    input px2777 ;
    input px2780 ;
    output px3304 ;
    output px3305 ;
    input px2841 ;
    input px2866 ;
    input px2821 ;
    input px2823 ;
    output px3359 ;
    input \p_key_samp(13)   ;
    output px3504 ;
    output px3723 ;
    output px3315 ;
    output px3316 ;
    output px3321 ;
    output px3322 ;
    input px2803 ;
    input px2810 ;
    input px2812 ;
    input \p_key_samp(6)   ;
    input px2801 ;
    input px2867 ;
    input px2827 ;
    input px2698 ;
    input px2702 ;
    input px2703 ;
    input \p_key_samp(61)   ;
    input px2733 ;
    input px2741 ;
    input px2723 ;
    input px2729 ;
    input px2711 ;
    input px2712 ;
    input px2764 ;
    input px2751 ;
    input \p_key_samp(10)   ;
    input \p_key_samp(46)   ;
    input px2680 ;
    input px2682 ;
    input px2683 ;
    input px2694 ;
    input \p_key_samp(21)   ;
    input \p_key_samp(12)   ;
    input \p_key_samp(5)   ;
    input \p_key_samp(7)   ;
    input px2765 ;
    input px2719 ;
    input px2709 ;
    input px2731 ;
    input \p_key_samp(49)   ;
    input px2642 ;
    input px2643 ;
    input px2644 ;
    input px2646 ;
    input px2618 ;
    input px2621 ;
    input px2622 ;
    input px2623 ;
    input \p_key_samp(39)   ;
    input \p_key_samp(47)   ;
    input \p_key_samp(28)   ;
    input px2654 ;
    input px2656 ;
    input px2658 ;
    input px2664 ;
    input \p_key_samp(23)   ;
    input px2630 ;
    input px2634 ;
    input px2637 ;
    input px2638 ;
    input \p_key_samp(22)   ;
    input \p_key_samp(54)   ;
    input \p_key_samp(37)   ;
    input px2668 ;
    input px2670 ;
    input px2669 ;
    input px2672 ;
    input px2605 ;
    input px2606 ;
    input px2607 ;
    input px2608 ;
    output px3007 ;
    input \p_key_samp(14)   ;
    input \p_key_samp(63)   ;
    input \p_key_samp(30)   ;
    input \p_key_samp(53)   ;
    input \p_key_samp(31)   ;
    input px2514 ;
    input px2507 ;
    input \p_key_samp(29)   ;
    input \p_key_samp(20)   ;
    output px3036 ;
    input \p_key_samp(62)   ;
    input \p_key_samp(38)   ;
    input \p_key_samp(55)   ;
    input px2497 ;
    input \p_key_samp(19)   ;
    input \p_key_samp(52)   ;
    output px3052 ;
    input \p_key_samp(59)   ;
    input \p_key_samp(34)   ;
    input \p_key_samp(2)   ;
    input \p_key_samp(17)   ;
    input \p_key_samp(26)   ;
    input px2585 ;
    input px2591 ;
    input px2587 ;
    input px2593 ;
    input \p_key_samp(51)   ;
    input \p_key_samp(3)   ;
    input \p_key_samp(33)   ;
    input \p_key_samp(9)   ;
    input px2628 ;
    input px2640 ;
    input px2678 ;
    input px2706 ;
    input \p_key_samp(27)   ;
    input \p_key_samp(35)   ;
    input \p_key_samp(58)   ;
    input px2570 ;
    input px2569 ;
    input px2566 ;
    input px2563 ;
    input \p_key_samp(36)   ;
    input px2573 ;
    input px2575 ;
    input px2579 ;
    input px2582 ;
    input \p_key_samp(18)   ;
    input px2601 ;
    input px2611 ;
    input px2613 ;
    input px2615 ;
    input \p_key_samp(41)   ;
    input px2551 ;
    input px2555 ;
    input px2557 ;
    input px2558 ;
    input \p_key_samp(60)   ;
    input \p_key_samp(25)   ;
    input \p_key_samp(42)   ;
    input \p_key_samp(1)   ;
    input \p_key_samp(11)   ;
    input px2528 ;
    input px2523 ;
    input px2522 ;
    input px2521 ;
    input \p_key_samp(57)   ;
    input px2537 ;
    input px2534 ;
    input px2533 ;
    input px2538 ;
    input \p_key_samp(43)   ;
    output px2708 ;
    output px2869 ;
    output px3058 ;
    output px3281 ;
    output px3503 ;
    output px2432 ;
    output px2707 ;
    output px2868 ;
    output px3057 ;
    output px3221 ;
    output px3222 ;
    output px2431 ;
    output px2430 ;
    output px2429 ;
    output px2576 ;
    output px2742 ;
    output px2891 ;
    output px3092 ;
    output px3093 ;
    output px2428 ;
    output px2588 ;
    output px2768 ;
    output px2941 ;
    output px3151 ;
    output px3152 ;
    output px2427 ;
    output px2426 ;
    output px2425 ;
    output px2592 ;
    output px2786 ;
    output px2945 ;
    output px3160 ;
    output px3161 ;
    output px2424 ;
    output px2641 ;
    output px2828 ;
    output px2953 ;
    output px3187 ;
    output px3202 ;
    output px2423 ;
    output px2422 ;
    output px2421 ;
    output px2420 ;
    output px2629 ;
    output px2802 ;
    output px3017 ;
    output px3170 ;
    output px3185 ;
    output px2419 ;
    output px2418 ;
    output px2556 ;
    output px2730 ;
    output px2899 ;
    output px3068 ;
    output px3069 ;
    output px2417 ;
    output px2602 ;
    output px2748 ;
    output px2914 ;
    output px3119 ;
    output px3120 ;
    output px2416 ;
    output px2415 ;
    output px2594 ;
    output px2772 ;
    output px2929 ;
    output px3138 ;
    output px3149 ;
    output px2414 ;
    output px2413 ;
    output px2614 ;
    output px2752 ;
    output px2909 ;
    output px3112 ;
    output px3113 ;
    output px2412 ;
    output px2586 ;
    output px2770 ;
    output px2943 ;
    output px3154 ;
    output px3155 ;
    output px2411 ;
    output px2410 ;
    output px2409 ;
    output px2552 ;
    output px2728 ;
    output px2895 ;
    output px3073 ;
    output px3074 ;
    output px2408 ;
    output px2574 ;
    output px2734 ;
    output px2885 ;
    output px3095 ;
    output px3096 ;
    output px2407 ;
    output px2406 ;
    output px2405 ;
    output px2612 ;
    output px2746 ;
    output px2907 ;
    output px3109 ;
    output px3110 ;
    output px2404 ;
    output px2403 ;
    output px2402 ;
    output px2679 ;
    output px2790 ;
    output px2985 ;
    output px3245 ;
    output px3280 ;
    output px2401 ;
    output px2671 ;
    output px2855 ;
    output px3010 ;
    output px3216 ;
    output px3217 ;
    output px2400 ;
    output px2639 ;
    output px2807 ;
    output px3022 ;
    output px3172 ;
    output px3173 ;
    output px2399 ;
    output px2665 ;
    output px2820 ;
    output px2973 ;
    output px3232 ;
    output px3233 ;
    output px2398 ;
    output px2766 ;
    output px2927 ;
    output px3136 ;
    output px3330 ;
    output px3349 ;
    output px2397 ;
    output px2396 ;
    output px2395 ;
    output px2394 ;
    output px2393 ;
    output px2392 ;
    output px2391 ;
    output px2390 ;
    output px2389 ;
    output px2720 ;
    output px2893 ;
    output px3060 ;
    output px3296 ;
    output px3311 ;
    output px2388 ;
    output px2647 ;
    output px2832 ;
    output px3054 ;
    output px3197 ;
    output px3198 ;
    output px2387 ;
    output px2655 ;
    output px2818 ;
    output px2970 ;
    output px3229 ;
    output px3230 ;
    output px2386 ;
    output px2695 ;
    output px2798 ;
    output px2997 ;
    output px3278 ;
    output px3279 ;
    output px2385 ;
    output px2710 ;
    output px2871 ;
    output px3077 ;
    output px3283 ;
    output px3294 ;
    output px2384 ;
    output px2508 ;
    output px2645 ;
    output px2836 ;
    output px3035 ;
    output px3191 ;
    output px3192 ;
    output px2383 ;
    output px2657 ;
    output px2822 ;
    output px2967 ;
    output px3226 ;
    output px3227 ;
    output px2382 ;
    output px2681 ;
    output px2795 ;
    output px2987 ;
    output px3261 ;
    output px3262 ;
    output px2381 ;
    output px2380 ;
    output px2379 ;
    output px2378 ;
    output px2377 ;
    output px2376 ;
    output px2375 ;
    output px2374 ;
    output px2373 ;
    output px2732 ;
    output px2881 ;
    output px3090 ;
    output px3313 ;
    output px3328 ;
    output px2372 ;
    output px2520 ;
    output px2673 ;
    output px2857 ;
    output px3006 ;
    output px3206 ;
    output px3207 ;
    output px2371 ;
    output px2498 ;
    output px2631 ;
    output px2811 ;
    output px3041 ;
    output px3183 ;
    output px3184 ;
    output px2370 ;
    output px2659 ;
    output px2824 ;
    output px2982 ;
    output px3235 ;
    output px3236 ;
    output px2369 ;
    input [63:0]p_nbus_data_in_int ;
    output [63:63]p_nbus_plaintext ;
    output \p_plaintext(37)   ;
    output \p_plaintext(39)   ;
    input p_reset_int ;
    input p_load_int ;
    input p_clk_int ;
    output \p_plaintext(63)   ;

    wire nx63157z22, nx63157z24, nx63157z26, nx63157z23, nx63157z21, nx63157z25, 
         nx63157z9, nx63157z8, nx63157z10, nx63157z6, nx63157z5, nx63157z7, 
         nx40221z8, nx40221z7, nx40221z6, nx40221z5, nx40221z4, nx40221z3, 
         nx39226z13, nx39226z12, nx39226z10, nx39226z8, nx63157z50, nx63157z49, 
         nx63157z48, nx63157z47, nx63157z46, nx63157z45, nx63157z14, nx63157z16, 
         nx63157z18, nx63157z15, nx63157z13, nx63157z34, nx63157z33, nx63157z32, 
         nx63157z31, nx63157z30, nx63157z29, nx63157z39, nx63157z42, nx63157z38, 
         nx63157z37, nx63157z40, nx63157z41, nx39226z14, nx39226z5, nx39226z18, 
         nx39226z3, nx39226z16, nx39226z6, nx63157z19, nx63157z11, nx63157z3, 
         nx63157z35, nx63157z43, nx63157z27, nx37232z12, nx37232z10, nx37232z8, 
         nx37232z7, nx37232z5, nx37232z3, nx34235z29, nx34235z27, nx34235z26, 
         nx34235z24, nx34235z23, nx34235z22, nx36228z12, nx36228z11, nx36228z9, 
         nx36228z7, nx36228z5, nx36228z3, nx34235z11, nx34235z19, nx34235z14, 
         nx34235z12, nx34235z16, nx34235z17, nx34235z35, nx34235z33, nx34235z36, 
         nx34235z38, nx34235z32, nx34235z39, nx29253z6, nx29253z9, nx29253z7, 
         nx29253z4, nx29253z5, nx29253z3, nx27254z12, nx27254z10, nx27254z8, 
         nx27254z6, nx27254z5, nx27254z3, nx15291z23, nx15291z22, nx15291z21, 
         nx15291z20, nx15291z17, nx15291z34, nx15291z33, nx15291z31, nx15291z30, 
         nx15291z28, nx15291z27, nx16286z4, nx16286z10, nx16286z5, nx16286z3, 
         nx16286z7, nx16286z8, nx16289z9, nx16289z6, nx16289z3, nx16289z8, 
         nx16289z4, nx34235z30, nx34235z20, nx34235z9, nx34235z7, nx34235z5, 
         nx34235z3, nx25263z10, nx25263z9, nx25263z7, nx25263z5, nx25263z4, 
         nx25263z3, nx15291z11, nx15291z10, nx15291z9, nx15291z7, nx15291z6, 
         nx15291z5, nx36230z10, nx36230z8, nx36230z4, nx36230z9, nx36230z2, 
         nx36230z6, nx37234z5, nx37234z8, nx37234z9, nx37234z4, nx37234z2, 
         nx37234z6, nx24265z32, nx24265z28, nx24265z34, nx24265z27, nx24265z29, 
         nx24265z30, nx24265z11, nx24265z10, nx24265z9, nx24265z8, nx24265z6, 
         nx24265z4, nx24265z24, nx24265z21, nx24265z22, nx24265z18, nx24265z19, 
         nx24265z17, nx13298z16, nx13298z19, nx13298z12, nx13298z17, nx13298z18, 
         nx13298z14, nx7313z11, nx7313z9, nx7313z8, nx7313z6, nx7313z5, nx7313z3, 
         nx15291z37, nx15291z35, nx15291z25, nx15291z15, nx15291z13, nx15291z3, 
         nx13298z20, nx13298z10, nx13298z8, nx13298z7, nx13298z6, nx13298z4, 
         nx13298z78, nx13298z77, nx13298z75, nx13298z74, nx13298z73, nx13298z71, 
         nx13298z51, nx13298z53, nx13298z49, nx13298z58, nx13298z55, nx13298z57, 
         nx13298z34, nx13298z32, nx13298z30, nx13298z28, nx13298z26, nx13298z24, 
         nx13298z68, nx13298z67, nx13298z66, nx13298z64, nx13298z63, nx13298z61, 
         nx7312z16, nx7312z15, nx7312z14, nx7312z13, nx7312z11, nx7312z10, 
         nx13298z44, nx13298z45, nx13298z38, nx13298z40, nx13298z42, nx13298z41, 
         nx24265z2, nx24265z36, nx24265z35, nx24265z25, nx24265z15, nx24265z13, 
         nx5318z7, nx5318z4, nx5318z8, nx5318z5, nx5318z3, nx5318z2, nx9305z9, 
         nx9305z8, nx9305z7, nx9305z6, nx9305z4, nx9305z2, nx337z7, nx337z5, 
         nx337z2, nx337z8, nx337z3, nx337z9, nx11304z9, nx11304z8, nx11304z7, 
         nx11304z5, nx11304z4, nx11304z2, nx4319z9, nx4319z8, nx4319z7, nx4319z6, 
         nx4319z4, nx4319z2, nx3326z9, nx3326z7, nx3326z6, nx3326z4, nx3326z3, 
         nx3326z2, nx7312z6, nx7312z20, nx7312z2, nx7312z4, nx7312z18, nx7312z8, 
         nx13298z69, nx13298z59, nx13298z47, nx13298z36, nx13298z22, nx13298z2, 
         nx16286z9, nx16286z6, nx35956z10, nx35956z9, nx35956z8, nx35956z7, 
         nx35956z5, nx35956z3, nx32966z10, nx32966z8, nx32966z6, nx32966z5, 
         nx32966z4, nx32966z3, nx12903z12, nx12903z11, nx12903z9, nx12903z10, 
         nx12903z5, nx12903z7, nx12903z59, nx12903z57, nx12903z56, nx12903z54, 
         nx12903z53, nx12903z52, nx63157z4, nx37234z3, nx12903z341, nx63157z20, 
         nx27254z11, nx27254z9, nx12903z47, nx12903z43, nx12903z40, nx12903z42, 
         nx12903z44, nx12903z45, nx12903z19, nx12903z18, nx12903z24, nx12903z25, 
         nx12903z23, nx12903z21, nx63157z12, nx12903z78, nx12903z76, nx12903z75, 
         nx12903z74, nx12903z73, nx12903z72, nx12903z37, nx12903z35, nx12903z34, 
         nx12903z33, nx12903z32, nx12903z30, nx15291z8, nx15291z12, nx37234z7, 
         nx12903z343, nx63157z28, nx38222z2, nx12903z50, nx12903z48, nx12903z38, 
         nx12903z28, nx12903z26, nx12903z16, nx16289z10, nx16289z7, nx37232z2, 
         nx63157z44, nx39226z2, nx27254z4, nx25263z6, nx36228z2, nx25263z8, 
         nx27254z7, nx63157z36, nx12903z149, nx12903z148, nx12903z146, 
         nx12903z144, nx12903z143, nx12903z142, nx34235z10, nx34235z31, 
         nx12903z92, nx12903z87, nx12903z91, nx12903z84, nx12903z86, nx12903z89, 
         nx34235z4, nx12903z114, nx12903z113, nx12903z112, nx12903z110, 
         nx12903z108, nx12903z106, nx34235z8, nx37232z11, nx36228z6, nx34235z21, 
         nx12903z162, nx12903z161, nx12903z159, nx12903z158, nx12903z157, 
         nx12903z156, nx15291z24, nx12903z98, nx12903z102, nx12903z96, 
         nx12903z95, nx12903z103, nx12903z100, nx13298z54, nx15291z18, nx34235z6, 
         nx28253z2, nx36228z8, nx15291z36, nx12903z270, nx37232z9, nx36228z10, 
         nx12903z80, nx12903z70, nx12903z68, nx12903z66, nx12903z64, nx12903z62, 
         nx15291z32, nx12903z124, nx12903z122, nx12903z120, nx12903z119, 
         nx12903z118, nx12903z117, nx15291z29, nx23267z2, nx63157z2, nx29253z2, 
         nx36228z4, nx15291z38, nx12903z283, nx34235z37, nx13298z13, nx12903z134, 
         nx37232z13, nx40221z2, nx34235z34, nx13298z15, nx12903z170, nx13298z76, 
         nx12903z130, nx39226z15, nx39226z4, nx24265z7, nx12903z293, nx27254z2, 
         nx12903z296, nx39226z7, nx24265z12, nx12903z299, nx39226z17, nx44209z2, 
         nx12903z82, nx12903z93, nx12903z115, nx12903z14, nx12903z60, 
         nx12903z104, nx34235z15, nx12903z172, nx12903z178, nx12903z174, 
         nx12903z180, nx12903z176, nx12903z182, nx7313z4, nx12903z190, 
         nx34235z13, nx12903z205, nx12903z203, nx12903z201, nx12903z199, 
         nx12903z197, nx12903z195, nx7313z10, nx12903z193, nx34235z18, 
         nx12903z154, nx12903z138, nx12903z140, nx12903z136, nx12903z150, 
         nx12903z152, nx41222z2, nx45210z2, nx13298z72, nx12903z186, nx37232z6, 
         nx36230z5, nx12903z351, nx37232z4, nx36230z3, nx12903z355, nx36230z11, 
         nx12903z165, nx11304z3, nx61487z3, nx13298z5, nx12903z265, nx13298z9, 
         nx12903z288, nx29253z8, nx12903z236, nx12903z234, nx12903z233, 
         nx12903z231, nx12903z230, nx12903z229, nx24265z20, nx12903z227, 
         nx29253z10, nx12903z250, nx12903z249, nx12903z248, nx12903z247, 
         nx12903z245, nx12903z243, nx24265z23, nx12903z241, nx12903z364, 
         nx12903z358, nx12903z361, nx12903z362, nx12903z359, nx12903z357, 
         nx12903z400, nx34235z28, nx12903z278, nx12903z276, nx12903z275, 
         nx12903z274, nx12903z273, nx12903z272, nx24265z33, nx12903z404, 
         nx13298z39, nx12903z395, nx13298z46, nx12903z410, nx11304z6, nx61487z6, 
         nx13298z62, nx12903z335, nx12903z366, nx12903z365, nx12903z354, 
         nx12903z350, nx13298z65, nx12903z347, nx12903z298, nx12903z292, 
         nx12903z295, nx7312z17, nx12903z429, nx7312z12, nx12903z435, 
         nx12903z340, nx12903z345, nx12903z342, nx24265z37, nx12903z441, 
         nx12903z399, nx12903z406, nx12903z403, nx24265z26, nx12903z446, 
         nx12903z240, nx12903z226, nx13298z50, nx12903z223, nx12903z169, 
         nx12903z164, nx12903z133, nx3326z5, nx12903z261, nx12903z192, 
         nx12903z189, nx13298z25, nx12903z307, nx12903z282, nx12903z269, 
         nx13298z29, nx12903z310, nx3326z8, nx12903z304, nx12903z6, nx12903z214, 
         nx9305z3, nx12903z460, nx9305z5, nx12903z457, nx12903z218, nx9305z10, 
         nx12903z258, nx12903z287, nx12903z264, nx7312z3, nx12903z322, nx7312z7, 
         nx12903z373, nx12903z8, nx12903z319, nx12903z129, nx12903z185, 
         nx13298z70, nx42825z31, nx13298z60, nx42825z37, nx12903z251, 
         nx12903z222, nx5318z6, nx12903z381, nx12903z309, nx12903z306, nx5318z9, 
         nx12903z388, nx35956z6, nx42825z54, nx35956z4, nx42825z47, nx12903z445, 
         nx12903z440, nx4319z5, nx12903z472, nx12903z331, nx12903z394, 
         nx12903z409, nx4319z3, nx12903z477, nx12903z346, nx12903z334, nx337z4, 
         nx12903z421, nx24265z31, nx34235z25, nx12903z434, nx12903z428, nx337z6, 
         nx12903z425, nx12903z327, nx12903z41, nx12903z417, nx12903z46, 
         nx12903z453, nx12903z387, nx12903z380, nx12903z31, nx42825z110, 
         nx12903z36, nx42825z113, nx42825z60, nx12903z79, nx42825z128, 
         nx12903z456, nx12903z464, nx12903z459, nx12903z455, nx12903z463, 
         nx12903z77, nx42825z132, nx12903z377, nx42825z50, nx12903z450, 
         nx12903z424, nx12903z437, nx12903z420, nx12903z22, nx42825z146, 
         nx61487z8, nx61487z2, nx61487z5, nx12903z20, nx42825z151, nx12903z476, 
         nx12903z475, nx12903z471, nx32966z7, nx42825z75, nx12903z303, 
         nx12903z257, nx12903z217, nx12903z260, nx32966z9, nx12903z252, 
         nx12903z372, nx12903z330, nx12903z326, nx12903z321, nx12903z55, 
         nx42825z15, nx12903z467, nx42825z36, nx42825z33, nx42825z30, nx12903z58, 
         nx42825z26, nx42825z59, nx42825z56, nx42825z43, nx42825z46, nx42825z53, 
         nx42825z49, nx42825z25, nx42825z22, nx42825z19, nx42825z18, nx42825z17, 
         nx42825z14, nx12903z376, nx12903z213, nx12903z318, nx42825z82, 
         nx42825z79, nx42825z74, nx42825z4, nx42825z112, nx42825z109, 
         nx42825z106, nx42825z103, nx42825z131, nx42825z127, nx42825z123, 
         nx42825z122, nx42825z150, nx42825z145, nx42825z153, nx42825z149, 
         nx12903z480, nx12903z466, nx12903z416, nx12903z452, nx42825z94, 
         nx42825z189, nx42825z185, nx12903z391, nx12903z2, nx42825z155, 
         nx42825z142, nx42825z119, nx42825z99, nx42825z162, nx42825z93, 
         nx42825z3, nx42825z237, nx42825z197, nx42825z221, nx42825z222, 
         nx43816z5, nx42825z238, nx42825z85, nx42825z71, nx42825z176, 
         nx42825z172, nx43816z9, nx42825z11, nx42825z40, nx42825z216, 
         nx42825z209, nx43816z21, nx43816z25, nx43816z7, nx43816z3, nx43816z8, 
         nx43816z4, nx43820z9, nx43816z22, nx43820z14, nx43820z4, nx43820z8, 
         nx43820z13, nx43820z11, nx43824z4, nx43824z8, nx43820z5, nx43824z19, 
         nx43824z15, nx43824z10, nx43824z7, nx43824z3, nx43824z16, nx44815z20, 
         nx44815z23, nx44815z22, nx44815z19, nx44815z18, nx44815z13, nx44815z9, 
         nx44815z3, nx44815z10, nx42825z167, nx42825z182, nx44819z5, nx44819z8, 
         nx44815z4, nx42825z67, nx42825z8, nx44819z15, nx44819z14, nx44819z10, 
         nx44819z7, nx44819z4, nx44819z3, nx44819z16, nx44819z11, nx42825z229, 
         nx42825z233, nx42825z206, nx42825z202, nx45810z10, nx42825z139, 
         nx42825z96, nx42825z249, nx42825z243, nx45810z19, nx45810z4, nx45810z5, 
         nx45810z18, nx45810z9, nx45810z12, nx45810z3, nx42825z198, nx45810z6, 
         nx42825z163, nx45810z13, nx43816z29, nx43816z32, nx45814z8, nx43816z11, 
         nx43816z16, nx45814z11, nx45814z10, nx45814z7, nx45814z6, nx45814z5, 
         nx45814z4, nx45814z3, nx42825z2, nx42826z2, nx42827z2, nx42825z235, 
         nx42825z152, nx12903z442, nx12903z235, nx42825z234, nx43815z2, 
         nx42825z245, nx42825z129, nx12903z336, nx12903z277, nx42825z244, 
         nx43816z2, nx43817z2, nx43818z2, nx43816z31, nx42825z83, nx12903z253, 
         nx12903z196, nx43816z30, nx43819z2, nx42825z10, nx12903z215, 
         nx12903z131, nx12903z94, nx42825z9, nx43820z2, nx43821z2, nx43822z2, 
         nx42825z251, nx42825z133, nx12903z348, nx12903z279, nx42825z250, 
         nx43823z2, nx42825z141, nx12903z454, nx12903z411, nx12903z246, 
         nx42825z140, nx43824z2, nx42825z169, nx42825z48, nx12903z266, 
         nx12903z175, nx42825z168, nx44812z2, nx44813z2, nx43816z18, nx42825z27, 
         nx12903z311, nx12903z139, nx43816z17, nx44814z2, nx44815z2, nx44816z2, 
         nx42825z208, nx42825z114, nx12903z436, nx12903z363, nx42825z207, 
         nx44817z2, nx44818z2, nx43816z34, nx42825z76, nx12903z224, nx12903z200, 
         nx43816z33, nx44819z2, nx44820z2, nx44821z2, nx43816z13, nx42825z16, 
         nx12903z308, nx12903z137, nx43816z12, nx45809z2, nx42825z69, 
         nx12903z320, nx12903z187, nx12903z61, nx42825z68, nx45810z2, nx45811z2, 
         nx45812z2, nx42825z231, nx42825z147, nx12903z447, nx12903z232, 
         nx42825z230, nx45813z2, nx42825z98, nx12903z418, nx12903z396, 
         nx12903z244, nx42825z97, nx45814z2, nx45815z2, nx42825z184, nx42825z55, 
         nx12903z289, nx12903z177, nx42825z183, nx45816z2, nx42825z204, 
         nx42825z111, nx12903z430, nx12903z360, nx42825z203, nx45817z2, 
         nx43816z24, nx43824z18, nx44819z13, nx42825z166, nx43816z6, nx42825z42, 
         nx12903z262, nx12903z171, nx12903z101, nx42825z41, nx43824z5, 
         nx42825z178, nx42825z38, nx12903z271, nx12903z121, nx42825z177, 
         nx44819z9, nx42825z73, nx12903z374, nx12903z194, nx12903z63, nx42825z72, 
         nx45814z9, nx42825z187, nx12903z382, nx12903z294, nx12903z27, 
         nx42825z186, nx43816z10, nx42825z13, nx12903z305, nx12903z135, 
         nx12903z99, nx42825z12, nx43824z9, nx42825z174, nx42825z32, nx12903z284, 
         nx12903z123, nx42825z173, nx44819z6, nx42825z87, nx12903z323, 
         nx12903z191, nx12903z65, nx42825z86, nx45814z12, nx42825z191, 
         nx12903z389, nx12903z300, nx12903z51, nx42825z190, nx42825z242, 
         nx43820z7, nx44815z12, nx45810z8, nx42825z226, nx44815z8, nx45810z17, 
         nx42825z5, nx12903z211, nx12903z126, nx12903z13, nx12903z4, nx12903z3, 
         nx43820z15, nx42825z144, nx12903z458, nx12903z352, nx12903z111, 
         nx42825z143, nx44815z21, nx42825z211, nx12903z473, nx12903z228, 
         nx12903z163, nx42825z210, nx45810z20, nx42825z121, nx12903z422, 
         nx12903z405, nx12903z145, nx42825z120, nx42825z95, nx12903z414, 
         nx12903z393, nx12903z344, nx12903z88, nx12903z392, nx43820z10, 
         nx42825z157, nx12903z461, nx12903z356, nx12903z107, nx42825z156, 
         nx44815z24, nx42825z218, nx12903z478, nx12903z242, nx12903z160, 
         nx42825z217, nx45810z11, nx42825z101, nx12903z426, nx12903z401, 
         nx12903z147, nx42825z100, nx42825z200, nx44819z20;
    wire [6:0]plaintext;
    wire \plaintext(7)  , \plaintext(8)  , \plaintext(9)  , \plaintext(10)  , 
         \plaintext(11)  , \plaintext(12)  , \plaintext(13)  , \plaintext(14)  , 
         \plaintext(15)  , \plaintext(16)  , \plaintext(17)  , \plaintext(18)  , 
         \plaintext(19)  , \plaintext(20)  , \plaintext(21)  , \plaintext(22)  , 
         \plaintext(23)  , \plaintext(24)  , \plaintext(25)  , \plaintext(26)  , 
         \plaintext(27)  , \plaintext(28)  , \plaintext(29)  , \plaintext(30)  , 
         \plaintext(31)  , \plaintext(32)  , \plaintext(33)  , \plaintext(34)  , 
         \plaintext(35)  , \plaintext(36)  , \plaintext(38)  , \plaintext(40)  , 
         \plaintext(41)  , \plaintext(42)  , \plaintext(43)  , \plaintext(44)  , 
         \plaintext(45)  , \plaintext(46)  , \plaintext(47)  , \plaintext(48)  , 
         \plaintext(49)  , \plaintext(50)  , \plaintext(51)  , \plaintext(52)  , 
         \plaintext(53)  , \plaintext(54)  , \plaintext(55)  , \plaintext(56)  , 
         \plaintext(57)  , \plaintext(58)  , \plaintext(59)  , \plaintext(60)  , 
         \plaintext(61)  , \plaintext(62)  ;



    FDRE \reg_data_out(63)  (.Q (\p_plaintext(63)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[0]), .R (p_reset_int)) ;
    FDRE \reg_data_out(62)  (.Q (\plaintext(62)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[1]), .R (p_reset_int)) ;
    FDRE \reg_data_out(61)  (.Q (\plaintext(61)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[2]), .R (p_reset_int)) ;
    FDRE \reg_data_out(60)  (.Q (\plaintext(60)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[3]), .R (p_reset_int)) ;
    FDRE \reg_data_out(59)  (.Q (\plaintext(59)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[4]), .R (p_reset_int)) ;
    FDRE \reg_data_out(58)  (.Q (\plaintext(58)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[5]), .R (p_reset_int)) ;
    FDRE \reg_data_out(57)  (.Q (\plaintext(57)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[6]), .R (p_reset_int)) ;
    FDRE \reg_data_out(56)  (.Q (\plaintext(56)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[7]), .R (p_reset_int)) ;
    FDRE \reg_data_out(55)  (.Q (\plaintext(55)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[8]), .R (p_reset_int)) ;
    FDRE \reg_data_out(54)  (.Q (\plaintext(54)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[9]), .R (p_reset_int)) ;
    FDRE \reg_data_out(53)  (.Q (\plaintext(53)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[10]), .R (p_reset_int)) ;
    FDRE \reg_data_out(52)  (.Q (\plaintext(52)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[11]), .R (p_reset_int)) ;
    FDRE \reg_data_out(51)  (.Q (\plaintext(51)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[12]), .R (p_reset_int)) ;
    FDRE \reg_data_out(50)  (.Q (\plaintext(50)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[13]), .R (p_reset_int)) ;
    FDRE \reg_data_out(49)  (.Q (\plaintext(49)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[14]), .R (p_reset_int)) ;
    FDRE \reg_data_out(48)  (.Q (\plaintext(48)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[15]), .R (p_reset_int)) ;
    FDRE \reg_data_out(47)  (.Q (\plaintext(47)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[16]), .R (p_reset_int)) ;
    FDRE \reg_data_out(46)  (.Q (\plaintext(46)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[17]), .R (p_reset_int)) ;
    FDRE \reg_data_out(45)  (.Q (\plaintext(45)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[18]), .R (p_reset_int)) ;
    FDRE \reg_data_out(44)  (.Q (\plaintext(44)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[19]), .R (p_reset_int)) ;
    FDRE \reg_data_out(43)  (.Q (\plaintext(43)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[20]), .R (p_reset_int)) ;
    FDRE \reg_data_out(42)  (.Q (\plaintext(42)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[21]), .R (p_reset_int)) ;
    FDRE \reg_data_out(41)  (.Q (\plaintext(41)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[22]), .R (p_reset_int)) ;
    FDRE \reg_data_out(40)  (.Q (\plaintext(40)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[23]), .R (p_reset_int)) ;
    FDRE \reg_data_out(39)  (.Q (\p_plaintext(39)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[24]), .R (p_reset_int)) ;
    FDRE \reg_data_out(38)  (.Q (\plaintext(38)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[25]), .R (p_reset_int)) ;
    FDRE \reg_data_out(37)  (.Q (\p_plaintext(37)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[26]), .R (p_reset_int)) ;
    FDRE \reg_data_out(36)  (.Q (\plaintext(36)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[27]), .R (p_reset_int)) ;
    FDRE \reg_data_out(35)  (.Q (\plaintext(35)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[28]), .R (p_reset_int)) ;
    FDRE \reg_data_out(34)  (.Q (\plaintext(34)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[29]), .R (p_reset_int)) ;
    FDRE \reg_data_out(33)  (.Q (\plaintext(33)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[30]), .R (p_reset_int)) ;
    FDRE \reg_data_out(32)  (.Q (\plaintext(32)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[31]), .R (p_reset_int)) ;
    FDRE \reg_data_out(31)  (.Q (\plaintext(31)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[32]), .R (p_reset_int)) ;
    FDRE \reg_data_out(30)  (.Q (\plaintext(30)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[33]), .R (p_reset_int)) ;
    FDRE \reg_data_out(29)  (.Q (\plaintext(29)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[34]), .R (p_reset_int)) ;
    FDRE \reg_data_out(28)  (.Q (\plaintext(28)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[35]), .R (p_reset_int)) ;
    FDRE \reg_data_out(27)  (.Q (\plaintext(27)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[36]), .R (p_reset_int)) ;
    FDRE \reg_data_out(26)  (.Q (\plaintext(26)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[37]), .R (p_reset_int)) ;
    FDRE \reg_data_out(25)  (.Q (\plaintext(25)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[38]), .R (p_reset_int)) ;
    FDRE \reg_data_out(24)  (.Q (\plaintext(24)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[39]), .R (p_reset_int)) ;
    FDRE \reg_data_out(23)  (.Q (\plaintext(23)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[40]), .R (p_reset_int)) ;
    FDRE \reg_data_out(22)  (.Q (\plaintext(22)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[41]), .R (p_reset_int)) ;
    FDRE \reg_data_out(21)  (.Q (\plaintext(21)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[42]), .R (p_reset_int)) ;
    FDRE \reg_data_out(20)  (.Q (\plaintext(20)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[43]), .R (p_reset_int)) ;
    FDRE \reg_data_out(19)  (.Q (\plaintext(19)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[44]), .R (p_reset_int)) ;
    FDRE \reg_data_out(18)  (.Q (\plaintext(18)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[45]), .R (p_reset_int)) ;
    FDRE \reg_data_out(17)  (.Q (\plaintext(17)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[46]), .R (p_reset_int)) ;
    FDRE \reg_data_out(16)  (.Q (\plaintext(16)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[47]), .R (p_reset_int)) ;
    FDRE \reg_data_out(15)  (.Q (\plaintext(15)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[48]), .R (p_reset_int)) ;
    FDRE \reg_data_out(14)  (.Q (\plaintext(14)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[49]), .R (p_reset_int)) ;
    FDRE \reg_data_out(13)  (.Q (\plaintext(13)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[50]), .R (p_reset_int)) ;
    FDRE \reg_data_out(12)  (.Q (\plaintext(12)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[51]), .R (p_reset_int)) ;
    FDRE \reg_data_out(11)  (.Q (\plaintext(11)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[52]), .R (p_reset_int)) ;
    FDRE \reg_data_out(10)  (.Q (\plaintext(10)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[53]), .R (p_reset_int)) ;
    FDRE \reg_data_out(9)  (.Q (\plaintext(9)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[54]), .R (p_reset_int)) ;
    FDRE \reg_data_out(8)  (.Q (\plaintext(8)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[55]), .R (p_reset_int)) ;
    FDRE \reg_data_out(7)  (.Q (\plaintext(7)  ), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[56]), .R (p_reset_int)) ;
    FDRE \reg_data_out(6)  (.Q (plaintext[0]), .C (p_clk_int), .CE (p_load_int)
         , .D (p_nbus_data_in_int[57]), .R (p_reset_int)) ;
    FDRE \reg_data_out(5)  (.Q (p_nbus_plaintext[63]), .C (p_clk_int), .CE (
         p_load_int), .D (p_nbus_data_in_int[58]), .R (p_reset_int)) ;
    FDRE \reg_data_out(4)  (.Q (plaintext[2]), .C (p_clk_int), .CE (p_load_int)
         , .D (p_nbus_data_in_int[59]), .R (p_reset_int)) ;
    FDRE \reg_data_out(3)  (.Q (plaintext[3]), .C (p_clk_int), .CE (p_load_int)
         , .D (p_nbus_data_in_int[60]), .R (p_reset_int)) ;
    FDRE \reg_data_out(2)  (.Q (plaintext[4]), .C (p_clk_int), .CE (p_load_int)
         , .D (p_nbus_data_in_int[61]), .R (p_reset_int)) ;
    FDRE \reg_data_out(1)  (.Q (plaintext[5]), .C (p_clk_int), .CE (p_load_int)
         , .D (p_nbus_data_in_int[62]), .R (p_reset_int)) ;
    FDRE \reg_data_out(0)  (.Q (plaintext[6]), .C (p_clk_int), .CE (p_load_int)
         , .D (p_nbus_data_in_int[63]), .R (p_reset_int)) ;
    LUT6 ix50796z39819 (.O (px2369), .I0 (px3236), .I1 (px3235), .I2 (px2982), .I3 (
         px2824), .I4 (px2659), .I5 (nx44819z20)) ;
         defparam ix50796z39819.INIT = 64'h9669699669969669;
    LUT6 ix49808z39819 (.O (px2370), .I0 (px3184), .I1 (px3183), .I2 (px3041), .I3 (
         px2811), .I4 (px2631), .I5 (px2498)) ;
         defparam ix49808z39819.INIT = 64'h9669699669969669;
    LUT6 ix49807z28344 (.O (px2371), .I0 (px3207), .I1 (px3206), .I2 (px3006), .I3 (
         px2857), .I4 (px2673), .I5 (px2520)) ;
         defparam ix49807z28344.INIT = 64'h6996966996696996;
    LUT6 ix49806z28344 (.O (px2372), .I0 (px3328), .I1 (px3313), .I2 (px3090), .I3 (
         px2881), .I4 (px2732), .I5 (nx42825z200)) ;
         defparam ix49806z28344.INIT = 64'h6996966996696996;
    LUT6 ix49805z39819 (.O (px2373), .I0 (nx42825z100), .I1 (nx12903z147), .I2 (
         nx12903z401), .I3 (nx12903z426), .I4 (nx42825z101), .I5 (nx45810z11)) ;
         defparam ix49805z39819.INIT = 64'h9669699669969669;
    LUT6 ix49804z28344 (.O (px2374), .I0 (nx42825z217), .I1 (nx12903z160), .I2 (
         nx12903z242), .I3 (nx12903z478), .I4 (nx42825z218), .I5 (nx44815z24)) ;
         defparam ix49804z28344.INIT = 64'h6996966996696996;
    LUT6 ix49803z39819 (.O (px2375), .I0 (nx42825z156), .I1 (nx12903z107), .I2 (
         nx12903z356), .I3 (nx12903z461), .I4 (nx42825z157), .I5 (nx43820z10)) ;
         defparam ix49803z39819.INIT = 64'h9669699669969669;
    LUT6 ix49802z28344 (.O (px2376), .I0 (nx12903z392), .I1 (nx12903z88), .I2 (
         nx12903z344), .I3 (nx12903z393), .I4 (nx12903z414), .I5 (nx42825z95)) ;
         defparam ix49802z28344.INIT = 64'h6996966996696996;
    LUT6 ix49801z39819 (.O (px2377), .I0 (nx42825z120), .I1 (nx12903z145), .I2 (
         nx12903z405), .I3 (nx12903z422), .I4 (nx42825z121), .I5 (nx45810z20)) ;
         defparam ix49801z39819.INIT = 64'h9669699669969669;
    LUT6 ix49800z39819 (.O (px2378), .I0 (nx42825z210), .I1 (nx12903z163), .I2 (
         nx12903z228), .I3 (nx12903z473), .I4 (nx42825z211), .I5 (nx44815z21)) ;
         defparam ix49800z39819.INIT = 64'h9669699669969669;
    LUT6 ix49799z28344 (.O (px2379), .I0 (nx42825z143), .I1 (nx12903z111), .I2 (
         nx12903z352), .I3 (nx12903z458), .I4 (nx42825z144), .I5 (nx43820z15)) ;
         defparam ix49799z28344.INIT = 64'h6996966996696996;
    LUT6 ix48811z39819 (.O (px2380), .I0 (nx12903z3), .I1 (nx12903z4), .I2 (
         nx12903z13), .I3 (nx12903z126), .I4 (nx12903z211), .I5 (nx42825z5)) ;
         defparam ix48811z39819.INIT = 64'h9669699669969669;
    LUT6 ix48810z39819 (.O (px2381), .I0 (px3262), .I1 (px3261), .I2 (px2987), .I3 (
         px2795), .I4 (px2681), .I5 (nx45810z17)) ;
         defparam ix48810z39819.INIT = 64'h9669699669969669;
    LUT6 ix48809z28344 (.O (px2382), .I0 (px3227), .I1 (px3226), .I2 (px2967), .I3 (
         px2822), .I4 (px2657), .I5 (nx44815z8)) ;
         defparam ix48809z28344.INIT = 64'h6996966996696996;
    LUT6 ix48808z39819 (.O (px2383), .I0 (px3192), .I1 (px3191), .I2 (px3035), .I3 (
         px2836), .I4 (px2645), .I5 (px2508)) ;
         defparam ix48808z39819.INIT = 64'h9669699669969669;
    LUT6 ix48807z28344 (.O (px2384), .I0 (px3294), .I1 (px3283), .I2 (px3077), .I3 (
         px2871), .I4 (px2710), .I5 (nx42825z226)) ;
         defparam ix48807z28344.INIT = 64'h6996966996696996;
    LUT6 ix48806z28344 (.O (px2385), .I0 (px3279), .I1 (px3278), .I2 (px2997), .I3 (
         px2798), .I4 (px2695), .I5 (nx45810z8)) ;
         defparam ix48806z28344.INIT = 64'h6996966996696996;
    LUT6 ix48805z39819 (.O (px2386), .I0 (px3230), .I1 (px3229), .I2 (px2970), .I3 (
         px2818), .I4 (px2655), .I5 (nx44815z12)) ;
         defparam ix48805z39819.INIT = 64'h9669699669969669;
    LUT6 ix48804z39819 (.O (px2387), .I0 (px3198), .I1 (px3197), .I2 (px3054), .I3 (
         px2832), .I4 (px2647), .I5 (nx43820z7)) ;
         defparam ix48804z39819.INIT = 64'h9669699669969669;
    LUT6 ix48803z39819 (.O (px2388), .I0 (px3311), .I1 (px3296), .I2 (px3060), .I3 (
         px2893), .I4 (px2720), .I5 (nx42825z242)) ;
         defparam ix48803z39819.INIT = 64'h9669699669969669;
    LUT6 ix48802z28344 (.O (px2389), .I0 (nx42825z190), .I1 (nx12903z51), .I2 (
         nx12903z300), .I3 (nx12903z389), .I4 (nx42825z191), .I5 (nx45814z12)) ;
         defparam ix48802z28344.INIT = 64'h6996966996696996;
    LUT6 ix47814z28344 (.O (px2390), .I0 (nx42825z86), .I1 (nx12903z65), .I2 (
         nx12903z191), .I3 (nx12903z323), .I4 (nx42825z87), .I5 (nx44819z6)) ;
         defparam ix47814z28344.INIT = 64'h6996966996696996;
    LUT6 ix47813z39819 (.O (px2391), .I0 (nx42825z173), .I1 (nx12903z123), .I2 (
         nx12903z284), .I3 (nx42825z32), .I4 (nx42825z174), .I5 (nx43824z9)) ;
         defparam ix47813z39819.INIT = 64'h9669699669969669;
    LUT6 ix47812z39819 (.O (px2392), .I0 (nx42825z12), .I1 (nx12903z99), .I2 (
         nx12903z135), .I3 (nx12903z305), .I4 (nx42825z13), .I5 (nx43816z10)) ;
         defparam ix47812z39819.INIT = 64'h9669699669969669;
    LUT6 ix47811z28344 (.O (px2393), .I0 (nx42825z186), .I1 (nx12903z27), .I2 (
         nx12903z294), .I3 (nx12903z382), .I4 (nx42825z187), .I5 (nx45814z9)) ;
         defparam ix47811z28344.INIT = 64'h6996966996696996;
    LUT6 ix47810z39819 (.O (px2394), .I0 (nx42825z72), .I1 (nx12903z63), .I2 (
         nx12903z194), .I3 (nx12903z374), .I4 (nx42825z73), .I5 (nx44819z9)) ;
         defparam ix47810z39819.INIT = 64'h9669699669969669;
    LUT6 ix47809z39819 (.O (px2395), .I0 (nx42825z177), .I1 (nx12903z121), .I2 (
         nx12903z271), .I3 (nx42825z38), .I4 (nx42825z178), .I5 (nx43824z5)) ;
         defparam ix47809z39819.INIT = 64'h9669699669969669;
    LUT6 ix47808z39819 (.O (px2396), .I0 (nx42825z41), .I1 (nx12903z101), .I2 (
         nx12903z171), .I3 (nx12903z262), .I4 (nx42825z42), .I5 (nx43816z6)) ;
         defparam ix47808z39819.INIT = 64'h9669699669969669;
    LUT6 ix47807z39819 (.O (px2397), .I0 (px3349), .I1 (px3330), .I2 (px3136), .I3 (
         px2927), .I4 (px2766), .I5 (nx42825z166)) ;
         defparam ix47807z39819.INIT = 64'h9669699669969669;
    LUT6 ix47806z39819 (.O (px2398), .I0 (px3233), .I1 (px3232), .I2 (px2973), .I3 (
         px2820), .I4 (px2665), .I5 (nx44819z13)) ;
         defparam ix47806z39819.INIT = 64'h9669699669969669;
    LUT6 ix47805z28344 (.O (px2399), .I0 (px3173), .I1 (px3172), .I2 (px3022), .I3 (
         px2807), .I4 (px2639), .I5 (nx43824z18)) ;
         defparam ix47805z28344.INIT = 64'h6996966996696996;
    LUT6 ix45818z28344 (.O (px2400), .I0 (px3217), .I1 (px3216), .I2 (px3010), .I3 (
         px2855), .I4 (px2671), .I5 (nx43816z24)) ;
         defparam ix45818z28344.INIT = 64'h6996966996696996;
    LUT6 ix45817z28344 (.O (px2401), .I0 (px3280), .I1 (px3245), .I2 (px2985), .I3 (
         px2790), .I4 (px2679), .I5 (nx45817z2)) ;
         defparam ix45817z28344.INIT = 64'h6996966996696996;
    LUT6 ix45816z39819 (.O (px2402), .I0 (nx42825z203), .I1 (nx12903z360), .I2 (
         nx12903z430), .I3 (nx42825z111), .I4 (nx42825z204), .I5 (nx45816z2)) ;
         defparam ix45816z39819.INIT = 64'h9669699669969669;
    LUT6 ix45815z28344 (.O (px2403), .I0 (nx42825z183), .I1 (nx12903z177), .I2 (
         nx12903z289), .I3 (nx42825z55), .I4 (nx42825z184), .I5 (nx45815z2)) ;
         defparam ix45815z28344.INIT = 64'h6996966996696996;
    LUT6 ix45814z28344 (.O (px2404), .I0 (px3110), .I1 (px3109), .I2 (px2907), .I3 (
         px2746), .I4 (px2612), .I5 (nx45814z2)) ;
         defparam ix45814z28344.INIT = 64'h6996966996696996;
    LUT6 ix45813z39819 (.O (px2405), .I0 (nx42825z97), .I1 (nx12903z244), .I2 (
         nx12903z396), .I3 (nx12903z418), .I4 (nx42825z98), .I5 (nx45813z2)) ;
         defparam ix45813z39819.INIT = 64'h9669699669969669;
    LUT6 ix45812z28344 (.O (px2406), .I0 (nx42825z230), .I1 (nx12903z232), .I2 (
         nx12903z447), .I3 (nx42825z147), .I4 (nx42825z231), .I5 (nx45812z2)) ;
         defparam ix45812z28344.INIT = 64'h6996966996696996;
    LUT6 ix45811z28344 (.O (px2407), .I0 (px3096), .I1 (px3095), .I2 (px2885), .I3 (
         px2734), .I4 (px2574), .I5 (nx45811z2)) ;
         defparam ix45811z28344.INIT = 64'h6996966996696996;
    LUT6 ix45810z39819 (.O (px2408), .I0 (px3074), .I1 (px3073), .I2 (px2895), .I3 (
         px2728), .I4 (px2552), .I5 (nx45810z2)) ;
         defparam ix45810z39819.INIT = 64'h9669699669969669;
    LUT6 ix45809z39819 (.O (px2409), .I0 (nx42825z68), .I1 (nx12903z61), .I2 (
         nx12903z187), .I3 (nx12903z320), .I4 (nx42825z69), .I5 (nx45809z2)) ;
         defparam ix45809z39819.INIT = 64'h9669699669969669;
    LUT6 ix44821z28344 (.O (px2410), .I0 (nx43816z12), .I1 (nx12903z137), .I2 (
         nx12903z308), .I3 (nx42825z16), .I4 (nx43816z13), .I5 (nx44821z2)) ;
         defparam ix44821z28344.INIT = 64'h6996966996696996;
    LUT6 ix44820z28344 (.O (px2411), .I0 (px3155), .I1 (px3154), .I2 (px2943), .I3 (
         px2770), .I4 (px2586), .I5 (nx44820z2)) ;
         defparam ix44820z28344.INIT = 64'h6996966996696996;
    LUT6 ix44819z28344 (.O (px2412), .I0 (px3113), .I1 (px3112), .I2 (px2909), .I3 (
         px2752), .I4 (px2614), .I5 (nx44819z2)) ;
         defparam ix44819z28344.INIT = 64'h6996966996696996;
    LUT6 ix44818z28344 (.O (px2413), .I0 (nx43816z33), .I1 (nx12903z200), .I2 (
         nx12903z224), .I3 (nx42825z76), .I4 (nx43816z34), .I5 (nx44818z2)) ;
         defparam ix44818z28344.INIT = 64'h6996966996696996;
    LUT6 ix44817z28344 (.O (px2414), .I0 (px3149), .I1 (px3138), .I2 (px2929), .I3 (
         px2772), .I4 (px2594), .I5 (nx44817z2)) ;
         defparam ix44817z28344.INIT = 64'h6996966996696996;
    LUT6 ix44816z28344 (.O (px2415), .I0 (nx42825z207), .I1 (nx12903z363), .I2 (
         nx12903z436), .I3 (nx42825z114), .I4 (nx42825z208), .I5 (nx44816z2)) ;
         defparam ix44816z28344.INIT = 64'h6996966996696996;
    LUT6 ix44815z28344 (.O (px2416), .I0 (px3120), .I1 (px3119), .I2 (px2914), .I3 (
         px2748), .I4 (px2602), .I5 (nx44815z2)) ;
         defparam ix44815z28344.INIT = 64'h6996966996696996;
    LUT6 ix44814z39819 (.O (px2417), .I0 (px3069), .I1 (px3068), .I2 (px2899), .I3 (
         px2730), .I4 (px2556), .I5 (nx44814z2)) ;
         defparam ix44814z39819.INIT = 64'h9669699669969669;
    LUT6 ix44813z28344 (.O (px2418), .I0 (nx43816z17), .I1 (nx12903z139), .I2 (
         nx12903z311), .I3 (nx42825z27), .I4 (nx43816z18), .I5 (nx44813z2)) ;
         defparam ix44813z28344.INIT = 64'h6996966996696996;
    LUT6 ix44812z28344 (.O (px2419), .I0 (px3185), .I1 (px3170), .I2 (px3017), .I3 (
         px2802), .I4 (px2629), .I5 (nx44812z2)) ;
         defparam ix44812z28344.INIT = 64'h6996966996696996;
    LUT6 ix43824z39819 (.O (px2420), .I0 (nx42825z168), .I1 (nx12903z175), .I2 (
         nx12903z266), .I3 (nx42825z48), .I4 (nx42825z169), .I5 (nx43824z2)) ;
         defparam ix43824z39819.INIT = 64'h9669699669969669;
    LUT6 ix43823z28344 (.O (px2421), .I0 (nx42825z140), .I1 (nx12903z246), .I2 (
         nx12903z411), .I3 (nx12903z454), .I4 (nx42825z141), .I5 (nx43823z2)) ;
         defparam ix43823z28344.INIT = 64'h6996966996696996;
    LUT6 ix43822z39819 (.O (px2422), .I0 (nx42825z250), .I1 (nx12903z279), .I2 (
         nx12903z348), .I3 (nx42825z133), .I4 (nx42825z251), .I5 (nx43822z2)) ;
         defparam ix43822z39819.INIT = 64'h9669699669969669;
    LUT6 ix43821z28344 (.O (px2423), .I0 (px3202), .I1 (px3187), .I2 (px2953), .I3 (
         px2828), .I4 (px2641), .I5 (nx43821z2)) ;
         defparam ix43821z28344.INIT = 64'h6996966996696996;
    LUT6 ix43820z39819 (.O (px2424), .I0 (px3161), .I1 (px3160), .I2 (px2945), .I3 (
         px2786), .I4 (px2592), .I5 (nx43820z2)) ;
         defparam ix43820z39819.INIT = 64'h9669699669969669;
    LUT6 ix43819z39819 (.O (px2425), .I0 (nx42825z9), .I1 (nx12903z94), .I2 (
         nx12903z131), .I3 (nx12903z215), .I4 (nx42825z10), .I5 (nx43819z2)) ;
         defparam ix43819z39819.INIT = 64'h9669699669969669;
    LUT6 ix43818z39819 (.O (px2426), .I0 (nx43816z30), .I1 (nx12903z196), .I2 (
         nx12903z253), .I3 (nx42825z83), .I4 (nx43816z31), .I5 (nx43818z2)) ;
         defparam ix43818z39819.INIT = 64'h9669699669969669;
    LUT6 ix43817z28344 (.O (px2427), .I0 (px3152), .I1 (px3151), .I2 (px2941), .I3 (
         px2768), .I4 (px2588), .I5 (nx43817z2)) ;
         defparam ix43817z28344.INIT = 64'h6996966996696996;
    LUT6 ix43816z39819 (.O (px2428), .I0 (px3093), .I1 (px3092), .I2 (px2891), .I3 (
         px2742), .I4 (px2576), .I5 (nx43816z2)) ;
         defparam ix43816z39819.INIT = 64'h9669699669969669;
    LUT6 ix43815z28344 (.O (px2429), .I0 (nx42825z244), .I1 (nx12903z277), .I2 (
         nx12903z336), .I3 (nx42825z129), .I4 (nx42825z245), .I5 (nx43815z2)) ;
         defparam ix43815z28344.INIT = 64'h6996966996696996;
    LUT6 ix42827z39819 (.O (px2430), .I0 (nx42825z234), .I1 (nx12903z235), .I2 (
         nx12903z442), .I3 (nx42825z152), .I4 (nx42825z235), .I5 (nx42827z2)) ;
         defparam ix42827z39819.INIT = 64'h9669699669969669;
    LUT6 ix42826z28344 (.O (px2431), .I0 (px3222), .I1 (px3221), .I2 (px3057), .I3 (
         px2868), .I4 (px2707), .I5 (nx42826z2)) ;
         defparam ix42826z28344.INIT = 64'h6996966996696996;
    LUT6 ix42825z28344 (.O (px2432), .I0 (px3503), .I1 (px3281), .I2 (px3058), .I3 (
         px2869), .I4 (px2708), .I5 (nx42825z2)) ;
         defparam ix42825z28344.INIT = 64'h6996966996696996;
    LUT6 ix45817z52308 (.O (nx45817z2), .I0 (nx45814z3), .I1 (nx45814z4), .I2 (
         nx45814z5), .I3 (nx45814z6), .I4 (nx45814z7), .I5 (nx45814z10)) ;
         defparam ix45817z52308.INIT = 64'hB64B2CC958A7C731;
    LUT6 ix45816z37254 (.O (nx45816z2), .I0 (nx45814z3), .I1 (nx45814z4), .I2 (
         nx45814z5), .I3 (nx45814z6), .I4 (nx45814z7), .I5 (nx45814z10)) ;
         defparam ix45816z37254.INIT = 64'h33E6C7583C998C63;
    LUT6 ix45815z28556 (.O (nx45815z2), .I0 (nx45814z3), .I1 (nx45814z4), .I2 (
         nx45814z5), .I3 (nx45814z6), .I4 (nx45814z7), .I5 (nx45814z10)) ;
         defparam ix45815z28556.INIT = 64'hA59356C6991E6A69;
    LUT6 ix45814z26205 (.O (nx45814z2), .I0 (nx45814z3), .I1 (nx45814z4), .I2 (
         nx45814z5), .I3 (nx45814z6), .I4 (nx45814z7), .I5 (nx45814z10)) ;
         defparam ix45814z26205.INIT = 64'hD38D9E640ED3613A;
    LUT6 ix45814z39828 (.O (nx45814z10), .I0 (\p_key_samp(43)  ), .I1 (
         nx45814z11), .I2 (nx12903z300), .I3 (nx12903z389), .I4 (nx42825z191), .I5 (
         nx45814z12)) ;
         defparam ix45814z39828.INIT = 64'h9669699669969669;
    LUT6 ix45814z36007 (.O (nx45814z12), .I0 (px2538), .I1 (px2533), .I2 (px2534
         ), .I3 (px2537), .I4 (nx43816z16), .I5 (nx43816z11)) ;
         defparam ix45814z36007.INIT = 64'hCA4434EF7186877A;
    LUT6 ix45814z28350 (.O (nx45814z7), .I0 (\p_key_samp(57)  ), .I1 (nx45814z8)
         , .I2 (nx12903z294), .I3 (nx12903z382), .I4 (nx42825z187), .I5 (
         nx45814z9)) ;
         defparam ix45814z28350.INIT = 64'h6996966996696996;
    LUT6 ix45814z57203 (.O (nx45814z9), .I0 (px2521), .I1 (px2522), .I2 (px2523)
         , .I3 (nx43816z32), .I4 (nx43816z29), .I5 (px2528)) ;
         defparam ix45814z57203.INIT = 64'hDB6C318629B3DA49;
    LUT6 ix45814z28349 (.O (nx45814z6), .I0 (\p_key_samp(11)  ), .I1 (nx45810z13
         ), .I2 (px2987), .I3 (px2795), .I4 (px2681), .I5 (nx45810z17)) ;
         defparam ix45814z28349.INIT = 64'h6996966996696996;
    LUT6 ix45814z39823 (.O (nx45814z5), .I0 (\p_key_samp(1)  ), .I1 (nx42825z163
         ), .I2 (px3136), .I3 (px2927), .I4 (px2766), .I5 (nx42825z166)) ;
         defparam ix45814z39823.INIT = 64'h9669699669969669;
    LUT6 ix45814z28347 (.O (nx45814z4), .I0 (\p_key_samp(42)  ), .I1 (nx45810z6)
         , .I2 (px2997), .I3 (px2798), .I4 (px2695), .I5 (nx45810z8)) ;
         defparam ix45814z28347.INIT = 64'h6996966996696996;
    LUT6 ix45814z39821 (.O (nx45814z3), .I0 (\p_key_samp(25)  ), .I1 (
         nx42825z198), .I2 (px3090), .I3 (px2881), .I4 (px2732), .I5 (
         nx42825z200)) ;
         defparam ix45814z39821.INIT = 64'h9669699669969669;
    LUT6 ix45813z26751 (.O (nx45813z2), .I0 (nx45810z3), .I1 (nx45810z12), .I2 (
         nx45810z9), .I3 (nx45810z18), .I4 (nx45810z5), .I5 (nx45810z4)) ;
         defparam ix45813z26751.INIT = 64'h63D49CA3B469635C;
    LUT6 ix45812z44139 (.O (nx45812z2), .I0 (nx45810z12), .I1 (nx45810z3), .I2 (
         nx45810z5), .I3 (nx45810z4), .I4 (nx45810z18), .I5 (nx45810z9)) ;
         defparam ix45812z44139.INIT = 64'h36C3C8B5393EA748;
    LUT6 ix45811z5997 (.O (nx45811z2), .I0 (nx45810z3), .I1 (nx45810z4), .I2 (
         nx45810z5), .I3 (nx45810z9), .I4 (nx45810z12), .I5 (nx45810z18)) ;
         defparam ix45811z5997.INIT = 64'h2B92D46D6DF6124A;
    LUT6 ix45810z19901 (.O (nx45810z2), .I0 (nx45810z3), .I1 (nx45810z4), .I2 (
         nx45810z5), .I3 (nx45810z9), .I4 (nx45810z12), .I5 (nx45810z18)) ;
         defparam ix45810z19901.INIT = 64'h1DDAE137A669489A;
    LUT6 ix45810z39836 (.O (nx45810z18), .I0 (\p_key_samp(60)  ), .I1 (
         nx45810z19), .I2 (nx12903z405), .I3 (nx12903z422), .I4 (nx42825z121), .I5 (
         nx45810z20)) ;
         defparam ix45810z39836.INIT = 64'h9669699669969669;
    LUT6 ix45810z23488 (.O (nx45810z20), .I0 (nx42825z243), .I1 (px2558), .I2 (
         px2557), .I3 (px2555), .I4 (nx42825z249), .I5 (px2551)) ;
         defparam ix45810z23488.INIT = 64'hE9061AF45AB5568B;
    LUT6 ix45810z28355 (.O (nx45810z12), .I0 (\p_key_samp(41)  ), .I1 (
         nx45810z13), .I2 (px2987), .I3 (px2795), .I4 (px2681), .I5 (nx45810z17)
         ) ;
         defparam ix45810z28355.INIT = 64'h6996966996696996;
    LUT6 ix45810z28812 (.O (nx45810z17), .I0 (nx42825z96), .I1 (px2615), .I2 (
         px2613), .I3 (px2611), .I4 (px2601), .I5 (nx42825z139)) ;
         defparam ix45810z28812.INIT = 64'h87692CD2B4A56B5A;
    LUT5 ix45810z28352 (.O (nx45810z9), .I0 (\p_key_samp(18)  ), .I1 (nx45810z10
         ), .I2 (nx12903z426), .I3 (nx42825z101), .I4 (nx45810z11)) ;
         defparam ix45810z28352.INIT = 32'h96696996;
    LUT6 ix45810z55477 (.O (nx45810z11), .I0 (px2582), .I1 (nx42825z202), .I2 (
         px2579), .I3 (nx42825z206), .I4 (px2575), .I5 (px2573)) ;
         defparam ix45810z55477.INIT = 64'h6B6624DA147BD389;
    LUT6 ix45810z28348 (.O (nx45810z5), .I0 (\p_key_samp(36)  ), .I1 (nx45810z6)
         , .I2 (px2997), .I3 (px2798), .I4 (px2695), .I5 (nx45810z8)) ;
         defparam ix45810z28348.INIT = 64'h6996966996696996;
    LUT6 ix45810z39827 (.O (nx45810z8), .I0 (nx42825z233), .I1 (nx42825z229), .I2 (
         px2563), .I3 (px2566), .I4 (px2569), .I5 (px2570)) ;
         defparam ix45810z39827.INIT = 64'h8DE3789CC31C966A;
    LUT6 ix45810z28347 (.O (nx45810z4), .I0 (\p_key_samp(58)  ), .I1 (nx44819z11
         ), .I2 (px2973), .I3 (px2820), .I4 (px2665), .I5 (nx44819z13)) ;
         defparam ix45810z28347.INIT = 64'h6996966996696996;
    LUT6 ix45810z28346 (.O (nx45810z3), .I0 (\p_key_samp(35)  ), .I1 (nx44819z16
         ), .I2 (px2982), .I3 (px2824), .I4 (px2659), .I5 (nx44819z20)) ;
         defparam ix45810z28346.INIT = 64'h6996966996696996;
    LUT6 ix45809z44219 (.O (nx45809z2), .I0 (nx44819z3), .I1 (nx44819z4), .I2 (
         nx44819z7), .I3 (nx44819z10), .I4 (nx44819z14), .I5 (nx44819z15)) ;
         defparam ix45809z44219.INIT = 64'h66A52778985BA798;
    LUT6 ix44821z23437 (.O (nx44821z2), .I0 (nx44819z4), .I1 (nx44819z15), .I2 (
         nx44819z3), .I3 (nx44819z7), .I4 (nx44819z10), .I5 (nx44819z14)) ;
         defparam ix44821z23437.INIT = 64'hD22DA75439C6566A;
    LUT6 ix44820z52030 (.O (nx44820z2), .I0 (nx44819z7), .I1 (nx44819z3), .I2 (
         nx44819z4), .I3 (nx44819z15), .I4 (nx44819z14), .I5 (nx44819z10)) ;
         defparam ix44820z52030.INIT = 64'h948B4BB46B3CC61B;
    LUT6 ix44819z54849 (.O (nx44819z2), .I0 (nx44819z3), .I1 (nx44819z4), .I2 (
         nx44819z7), .I3 (nx44819z10), .I4 (nx44819z14), .I5 (nx44819z15)) ;
         defparam ix44819z54849.INIT = 64'h361E6DA11DE1D11E;
    LUT6 ix44819z28358 (.O (nx44819z15), .I0 (\p_key_samp(27)  ), .I1 (
         nx44819z16), .I2 (px2982), .I3 (px2824), .I4 (px2659), .I5 (nx44819z20)
         ) ;
         defparam ix44819z28358.INIT = 64'h6996966996696996;
    LUT6 ix44819z19166 (.O (nx44819z20), .I0 (px2706), .I1 (px2678), .I2 (
         nx42825z8), .I3 (nx42825z67), .I4 (px2640), .I5 (px2628)) ;
         defparam ix44819z19166.INIT = 64'hEB0559E3965A45A9;
    LUT6 ix44819z28357 (.O (nx44819z14), .I0 (\p_key_samp(9)  ), .I1 (nx44815z4)
         , .I2 (px2967), .I3 (px2822), .I4 (px2657), .I5 (nx44815z8)) ;
         defparam ix44819z28357.INIT = 64'h6996966996696996;
    LUT6 ix44819z28353 (.O (nx44819z10), .I0 (\p_key_samp(33)  ), .I1 (
         nx44819z11), .I2 (px2973), .I3 (px2820), .I4 (px2665), .I5 (nx44819z13)
         ) ;
         defparam ix44819z28353.INIT = 64'h6996966996696996;
    LUT6 ix44819z36775 (.O (nx44819z13), .I0 (px2533), .I1 (px2534), .I2 (px2537
         ), .I3 (px2538), .I4 (nx43816z16), .I5 (nx43816z11)) ;
         defparam ix44819z36775.INIT = 64'hD33C6986A5C38A79;
    LUT6 ix44819z28350 (.O (nx44819z7), .I0 (\p_key_samp(3)  ), .I1 (nx44819z8)
         , .I2 (nx12903z194), .I3 (nx12903z374), .I4 (nx42825z73), .I5 (
         nx44819z9)) ;
         defparam ix44819z28350.INIT = 64'h6996966996696996;
    LUT6 ix44819z28113 (.O (nx44819z9), .I0 (px2528), .I1 (nx43816z29), .I2 (
         nx43816z32), .I3 (px2523), .I4 (px2522), .I5 (px2521)) ;
         defparam ix44819z28113.INIT = 64'hCC96A53197D868A7;
    LUT6 ix44819z28347 (.O (nx44819z4), .I0 (\p_key_samp(51)  ), .I1 (nx44819z5)
         , .I2 (nx12903z191), .I3 (nx12903z323), .I4 (nx42825z87), .I5 (
         nx44819z6)) ;
         defparam ix44819z28347.INIT = 64'h6996966996696996;
    LUT6 ix44819z15741 (.O (nx44819z6), .I0 (px2593), .I1 (px2587), .I2 (px2591)
         , .I3 (nx42825z182), .I4 (px2585), .I5 (nx42825z167)) ;
         defparam ix44819z15741.INIT = 64'h2C5587E9DAA53856;
    LUT6 ix44819z39821 (.O (nx44819z3), .I0 (\p_key_samp(26)  ), .I1 (nx44815z10
         ), .I2 (px2970), .I3 (px2818), .I4 (px2655), .I5 (nx44815z12)) ;
         defparam ix44819z39821.INIT = 64'h9669699669969669;
    LUT6 ix44818z52891 (.O (nx44818z2), .I0 (nx44815z3), .I1 (nx44815z9), .I2 (
         nx44815z13), .I3 (nx44815z18), .I4 (nx44815z19), .I5 (nx44815z22)) ;
         defparam ix44818z52891.INIT = 64'h1E6D51277689C978;
    LUT6 ix44817z43663 (.O (nx44817z2), .I0 (nx44815z3), .I1 (nx44815z9), .I2 (
         nx44815z13), .I3 (nx44815z18), .I4 (nx44815z19), .I5 (nx44815z22)) ;
         defparam ix44817z43663.INIT = 64'h79070AF1D61EA56C;
    LUT6 ix44816z16073 (.O (nx44816z2), .I0 (nx44815z13), .I1 (nx44815z3), .I2 (
         nx44815z19), .I3 (nx44815z18), .I4 (nx44815z9), .I5 (nx44815z22)) ;
         defparam ix44816z16073.INIT = 64'hC5365AC996C939A6;
    LUT6 ix44815z36856 (.O (nx44815z2), .I0 (nx44815z3), .I1 (nx44815z9), .I2 (
         nx44815z13), .I3 (nx44815z18), .I4 (nx44815z19), .I5 (nx44815z22)) ;
         defparam ix44815z36856.INIT = 64'hE34B69B21E688AD5;
    LUT6 ix44815z39840 (.O (nx44815z22), .I0 (\p_key_samp(17)  ), .I1 (
         nx44815z23), .I2 (nx12903z242), .I3 (nx12903z478), .I4 (nx42825z218), .I5 (
         nx44815z24)) ;
         defparam ix44815z39840.INIT = 64'h9669699669969669;
    LUT6 ix44815z15107 (.O (nx44815z24), .I0 (nx42825z96), .I1 (nx42825z139), .I2 (
         px2611), .I3 (px2613), .I4 (px2615), .I5 (px2601)) ;
         defparam ix44815z15107.INIT = 64'hCA5AA599363C35CA;
    LUT6 ix44815z28362 (.O (nx44815z19), .I0 (\p_key_samp(2)  ), .I1 (nx44815z20
         ), .I2 (nx12903z228), .I3 (nx12903z473), .I4 (nx42825z211), .I5 (
         nx44815z21)) ;
         defparam ix44815z28362.INIT = 64'h6996966996696996;
    LUT6 ix44815z44690 (.O (nx44815z21), .I0 (px2570), .I1 (px2569), .I2 (
         nx42825z229), .I3 (px2566), .I4 (nx42825z233), .I5 (px2563)) ;
         defparam ix44815z44690.INIT = 64'h47C9A9636C36A95C;
    LUT6 ix44815z39836 (.O (nx44815z18), .I0 (\p_key_samp(34)  ), .I1 (
         nx43824z16), .I2 (px3022), .I3 (px2807), .I4 (px2639), .I5 (nx43824z18)
         ) ;
         defparam ix44815z39836.INIT = 64'h9669699669969669;
    LUT6 ix44815z39831 (.O (nx44815z13), .I0 (\p_key_samp(59)  ), .I1 (px3052), 
         .I2 (px3041), .I3 (px2811), .I4 (px2631), .I5 (px2498)) ;
         defparam ix44815z39831.INIT = 64'h9669699669969669;
    LUT6 ix44815z39827 (.O (nx44815z9), .I0 (\p_key_samp(52)  ), .I1 (nx44815z10
         ), .I2 (px2970), .I3 (px2818), .I4 (px2655), .I5 (nx44815z12)) ;
         defparam ix44815z39827.INIT = 64'h9669699669969669;
    LUT6 ix44815z14745 (.O (nx44815z12), .I0 (nx42825z243), .I1 (px2558), .I2 (
         px2557), .I3 (px2555), .I4 (nx42825z249), .I5 (px2551)) ;
         defparam ix44815z14745.INIT = 64'h9B49C3B5C693346C;
    LUT6 ix44815z28346 (.O (nx44815z3), .I0 (\p_key_samp(19)  ), .I1 (nx44815z4)
         , .I2 (px2967), .I3 (px2822), .I4 (px2657), .I5 (nx44815z8)) ;
         defparam ix44815z28346.INIT = 64'h6996966996696996;
    LUT6 ix44815z40917 (.O (nx44815z8), .I0 (nx42825z202), .I1 (nx42825z206), .I2 (
         px2582), .I3 (px2579), .I4 (px2573), .I5 (px2575)) ;
         defparam ix44815z40917.INIT = 64'h295AC617C7639AAC;
    LUT6 ix44814z59064 (.O (nx44814z2), .I0 (nx43824z3), .I1 (px2497), .I2 (
         nx43824z7), .I3 (nx43824z10), .I4 (nx43824z15), .I5 (nx43824z19)) ;
         defparam ix44814z59064.INIT = 64'h95682AF27C8BE195;
    LUT6 ix44813z35961 (.O (nx44813z2), .I0 (nx43824z3), .I1 (px2497), .I2 (
         nx43824z7), .I3 (nx43824z10), .I4 (nx43824z15), .I5 (nx43824z19)) ;
         defparam ix44813z35961.INIT = 64'h56A1B9CBE01D8756;
    LUT6 ix44812z51638 (.O (nx44812z2), .I0 (px2497), .I1 (nx43824z10), .I2 (
         nx43824z3), .I3 (nx43824z7), .I4 (nx43824z15), .I5 (nx43824z19)) ;
         defparam ix44812z51638.INIT = 64'hAD67923C7AC1C493;
    LUT6 ix43824z54881 (.O (nx43824z2), .I0 (nx43824z3), .I1 (px2497), .I2 (
         nx43824z7), .I3 (nx43824z10), .I4 (nx43824z15), .I5 (nx43824z19)) ;
         defparam ix43824z54881.INIT = 64'h4F5416A9A987D13E;
    LUT6 ix43824z28361 (.O (nx43824z19), .I0 (\p_key_samp(55)  ), .I1 (nx43820z5
         ), .I2 (px3054), .I3 (px2832), .I4 (px2647), .I5 (nx43820z7)) ;
         defparam ix43824z28361.INIT = 64'h6996966996696996;
    LUT6 ix43824z39832 (.O (nx43824z15), .I0 (\p_key_samp(38)  ), .I1 (
         nx43824z16), .I2 (px3022), .I3 (px2807), .I4 (px2639), .I5 (nx43824z18)
         ) ;
         defparam ix43824z39832.INIT = 64'h9669699669969669;
    LUT6 ix43824z39118 (.O (nx43824z18), .I0 (nx43816z11), .I1 (px2538), .I2 (
         px2537), .I3 (nx43816z16), .I4 (px2534), .I5 (px2533)) ;
         defparam ix43824z39118.INIT = 64'h9B3CE8634669939C;
    LUT6 ix43824z28352 (.O (nx43824z10), .I0 (\p_key_samp(62)  ), .I1 (px3036), 
         .I2 (px3035), .I3 (px2836), .I4 (px2645), .I5 (px2508)) ;
         defparam ix43824z28352.INIT = 64'h6996966996696996;
    LUT6 ix43824z39824 (.O (nx43824z7), .I0 (\p_key_samp(20)  ), .I1 (nx43824z8)
         , .I2 (nx12903z284), .I3 (nx42825z32), .I4 (nx42825z174), .I5 (
         nx43824z9)) ;
         defparam ix43824z39824.INIT = 64'h9669699669969669;
    LUT6 ix43824z20167 (.O (nx43824z9), .I0 (nx42825z67), .I1 (px2706), .I2 (
         px2640), .I3 (px2678), .I4 (nx42825z8), .I5 (px2628)) ;
         defparam ix43824z20167.INIT = 64'h611EBC616EB1499E;
    LUT6 ix44815z16729 (.O (px2498), .I0 (px2523), .I1 (px2528), .I2 (nx43816z29
         ), .I3 (px2522), .I4 (px2521), .I5 (nx43816z32)) ;
         defparam ix44815z16729.INIT = 64'h671ACB84897D3C27;
    LUT6 ix43824z28346 (.O (nx43824z3), .I0 (\p_key_samp(29)  ), .I1 (nx43824z4)
         , .I2 (nx12903z271), .I3 (nx42825z38), .I4 (nx42825z178), .I5 (
         nx43824z5)) ;
         defparam ix43824z28346.INIT = 64'h6996966996696996;
    LUT6 ix43824z20112 (.O (nx43824z5), .I0 (nx42825z243), .I1 (px2558), .I2 (
         px2557), .I3 (px2555), .I4 (nx42825z249), .I5 (px2551)) ;
         defparam ix43824z20112.INIT = 64'h3C2D63D2DA69496A;
    LUT6 ix43823z39067 (.O (nx43823z2), .I0 (nx43820z11), .I1 (nx43820z13), .I2 (
         nx43820z8), .I3 (px2507), .I4 (nx43820z4), .I5 (px2514)) ;
         defparam ix43823z39067.INIT = 64'hB958CC874EA59378;
    LUT6 ix43822z12533 (.O (nx43822z2), .I0 (px2514), .I1 (nx43820z11), .I2 (
         nx43820z4), .I3 (nx43820z8), .I4 (nx43820z13), .I5 (px2507)) ;
         defparam ix43822z12533.INIT = 64'h7740D62C5CA72BD2;
    LUT6 ix43821z27580 (.O (nx43821z2), .I0 (px2514), .I1 (nx43820z4), .I2 (
         nx43820z8), .I3 (nx43820z11), .I4 (px2507), .I5 (nx43820z13)) ;
         defparam ix43821z27580.INIT = 64'h2D52D14E69B66699;
    LUT6 ix43820z52427 (.O (nx43820z2), .I0 (px2514), .I1 (nx43820z4), .I2 (
         nx43820z8), .I3 (nx43820z11), .I4 (px2507), .I5 (nx43820z13)) ;
         defparam ix43820z52427.INIT = 64'hC63938D6395AC7A8;
    LUT6 ix43820z28354 (.O (nx43820z13), .I0 (\p_key_samp(31)  ), .I1 (
         nx43820z14), .I2 (nx12903z352), .I3 (nx12903z458), .I4 (nx42825z144), .I5 (
         nx43820z15)) ;
         defparam ix43820z28354.INIT = 64'h6996966996696996;
    LUT6 ix43820z5007 (.O (nx43820z15), .I0 (px2570), .I1 (px2569), .I2 (
         nx42825z229), .I3 (px2566), .I4 (nx42825z233), .I5 (px2563)) ;
         defparam ix43820z5007.INIT = 64'hA49379E4799E0E61;
    LUT6 ix43824z52569 (.O (px2508), .I0 (nx42825z167), .I1 (px2593), .I2 (
         px2591), .I3 (nx42825z182), .I4 (px2587), .I5 (px2585)) ;
         defparam ix43824z52569.INIT = 64'hEB68129797D4C82B;
    LUT6 ix43820z28353 (.O (nx43820z11), .I0 (\p_key_samp(53)  ), .I1 (
         nx43816z22), .I2 (px3010), .I3 (px2855), .I4 (px2671), .I5 (nx43816z24)
         ) ;
         defparam ix43820z28353.INIT = 64'h6996966996696996;
    LUT6 ix43820z39825 (.O (nx43820z8), .I0 (\p_key_samp(30)  ), .I1 (nx43820z9)
         , .I2 (nx12903z356), .I3 (nx12903z461), .I4 (nx42825z157), .I5 (
         nx43820z10)) ;
         defparam ix43820z39825.INIT = 64'h9669699669969669;
    LUT6 ix43820z44047 (.O (nx43820z10), .I0 (nx42825z206), .I1 (nx42825z202), .I2 (
         px2582), .I3 (px2579), .I4 (px2575), .I5 (px2573)) ;
         defparam ix43820z44047.INIT = 64'hE86553393C92A6E5;
    LUT6 ix43820z28346 (.O (nx43820z4), .I0 (\p_key_samp(63)  ), .I1 (nx43820z5)
         , .I2 (px3054), .I3 (px2832), .I4 (px2647), .I5 (nx43820z7)) ;
         defparam ix43820z28346.INIT = 64'h6996966996696996;
    LUT6 ix43820z24237 (.O (nx43820z7), .I0 (nx42825z96), .I1 (px2615), .I2 (
         px2613), .I3 (px2611), .I4 (px2601), .I5 (nx42825z139)) ;
         defparam ix43820z24237.INIT = 64'h9AC365B9663C5986;
    LUT6 ix43819z24268 (.O (nx43819z2), .I0 (nx43816z4), .I1 (nx43816z8), .I2 (
         nx43816z3), .I3 (nx43816z7), .I4 (nx43816z25), .I5 (nx43816z21)) ;
         defparam ix43819z24268.INIT = 64'hCC63C3A53A5559A9;
    LUT6 ix43818z17021 (.O (nx43818z2), .I0 (nx43816z4), .I1 (nx43816z25), .I2 (
         nx43816z3), .I3 (nx43816z7), .I4 (nx43816z21), .I5 (nx43816z8)) ;
         defparam ix43818z17021.INIT = 64'hCD3253A896C53D5A;
    LUT6 ix43817z43897 (.O (nx43817z2), .I0 (nx43816z3), .I1 (nx43816z4), .I2 (
         nx43816z7), .I3 (nx43816z8), .I4 (nx43816z21), .I5 (nx43816z25)) ;
         defparam ix43817z43897.INIT = 64'h995A66697929A656;
    LUT6 ix43816z51853 (.O (nx43816z2), .I0 (nx43816z3), .I1 (nx43816z4), .I2 (
         nx43816z7), .I3 (nx43816z8), .I4 (nx43816z21), .I5 (nx43816z25)) ;
         defparam ix43816z51853.INIT = 64'h693C3AC53E91C56A;
    LUT6 ix43816z28364 (.O (nx43816z25), .I0 (\p_key_samp(14)  ), .I1 (px3007), 
         .I2 (px3006), .I3 (px2857), .I4 (px2673), .I5 (px2520)) ;
         defparam ix43816z28364.INIT = 64'h6996966996696996;
    LUT6 ix43816z27606 (.O (px2520), .I0 (px2528), .I1 (nx43816z29), .I2 (
         nx43816z32), .I3 (px2523), .I4 (px2522), .I5 (px2521)) ;
         defparam ix43816z27606.INIT = 64'h4FF8D027B844669E;
    LUT6 ix43816z28370 (.O (nx43816z32), .I0 (\p_key_samp(53)  ), .I1 (
         nx43816z33), .I2 (nx12903z200), .I3 (nx12903z224), .I4 (nx42825z76), .I5 (
         nx43816z34)) ;
         defparam ix43816z28370.INIT = 64'h6996966996696996;
    LUT6 ix43816z27416 (.O (nx43816z34), .I0 (nx42825z209), .I1 (px2608), .I2 (
         px2607), .I3 (px2606), .I4 (px2605), .I5 (nx42825z216)) ;
         defparam ix43816z27416.INIT = 64'hEDA6834C389665DA;
    LUT6 ix43816z39842 (.O (nx43816z29), .I0 (\p_key_samp(14)  ), .I1 (
         nx43816z30), .I2 (nx12903z196), .I3 (nx12903z253), .I4 (nx42825z83), .I5 (
         nx43816z31)) ;
         defparam ix43816z39842.INIT = 64'h9669699669969669;
    LUT6 ix43816z24551 (.O (nx43816z31), .I0 (nx42825z40), .I1 (px2672), .I2 (
         px2669), .I3 (px2670), .I4 (nx42825z11), .I5 (px2668)) ;
         defparam ix43816z24551.INIT = 64'h3AECE39645135AAC;
    LUT6 ix43816z28360 (.O (nx43816z21), .I0 (\p_key_samp(37)  ), .I1 (
         nx43816z22), .I2 (px3010), .I3 (px2855), .I4 (px2671), .I5 (nx43816z24)
         ) ;
         defparam ix43816z28360.INIT = 64'h6996966996696996;
    LUT6 ix43816z18671 (.O (nx43816z24), .I0 (px2640), .I1 (px2678), .I2 (
         nx42825z67), .I3 (px2706), .I4 (nx42825z8), .I5 (px2628)) ;
         defparam ix43816z18671.INIT = 64'h36C89525ADD643BA;
    LUT6 ix43816z39826 (.O (nx43816z8), .I0 (\p_key_samp(54)  ), .I1 (nx43816z9)
         , .I2 (nx12903z135), .I3 (nx12903z305), .I4 (nx42825z13), .I5 (
         nx43816z10)) ;
         defparam ix43816z39826.INIT = 64'h9669699669969669;
    LUT6 ix43816z56144 (.O (nx43816z10), .I0 (nx43816z11), .I1 (px2538), .I2 (
         px2537), .I3 (nx43816z16), .I4 (px2534), .I5 (px2533)) ;
         defparam ix43816z56144.INIT = 64'hC7262ADA38CBD625;
    LUT6 ix43816z28357 (.O (nx43816z16), .I0 (\p_key_samp(22)  ), .I1 (
         nx43816z17), .I2 (nx12903z139), .I3 (nx12903z311), .I4 (nx42825z27), .I5 (
         nx43816z18)) ;
         defparam ix43816z28357.INIT = 64'h6996966996696996;
    LUT6 ix43816z15224 (.O (nx43816z18), .I0 (px2638), .I1 (px2637), .I2 (
         nx42825z172), .I3 (px2634), .I4 (nx42825z176), .I5 (px2630)) ;
         defparam ix43816z15224.INIT = 64'hC235B5695CA93647;
    LUT6 ix43816z28354 (.O (nx43816z11), .I0 (\p_key_samp(23)  ), .I1 (
         nx43816z12), .I2 (nx12903z137), .I3 (nx12903z308), .I4 (nx42825z16), .I5 (
         nx43816z13)) ;
         defparam ix43816z28354.INIT = 64'h6996966996696996;
    LUT6 ix43816z30618 (.O (nx43816z13), .I0 (px2664), .I1 (nx42825z71), .I2 (
         nx42825z85), .I3 (px2658), .I4 (px2656), .I5 (px2654)) ;
         defparam ix43816z30618.INIT = 64'h72C99C966987726C;
    LUT6 ix43816z39825 (.O (nx43816z7), .I0 (\p_key_samp(28)  ), .I1 (
         nx42825z238), .I2 (px3060), .I3 (px2893), .I4 (px2720), .I5 (
         nx42825z242)) ;
         defparam ix43816z39825.INIT = 64'h9669699669969669;
    LUT6 ix43816z28347 (.O (nx43816z4), .I0 (\p_key_samp(47)  ), .I1 (
         nx12903z171), .I2 (nx43816z5), .I3 (nx12903z262), .I4 (nx42825z42), .I5 (
         nx43816z6)) ;
         defparam ix43816z28347.INIT = 64'h6996966996696996;
    LUT6 ix43816z9224 (.O (nx43816z6), .I0 (px2593), .I1 (nx42825z167), .I2 (
         px2591), .I3 (nx42825z182), .I4 (px2585), .I5 (px2587)) ;
         defparam ix43816z9224.INIT = 64'h9761D21E613E1EE1;
    LUT6 ix43816z28346 (.O (nx43816z3), .I0 (\p_key_samp(23)  ), .I1 (
         nx42825z222), .I2 (px3077), .I3 (px2871), .I4 (px2710), .I5 (
         nx42825z226)) ;
         defparam ix43816z28346.INIT = 64'h6996966996696996;
    LUT6 ix43815z39073 (.O (nx43815z2), .I0 (nx42825z221), .I1 (nx42825z197), .I2 (
         nx42825z237), .I3 (nx42825z3), .I4 (nx42825z93), .I5 (nx42825z162)) ;
         defparam ix43815z39073.INIT = 64'h167AEC8629C4937E;
    LUT6 ix42827z22479 (.O (nx42827z2), .I0 (nx42825z3), .I1 (nx42825z93), .I2 (
         nx42825z162), .I3 (nx42825z197), .I4 (nx42825z221), .I5 (nx42825z237)
         ) ;
         defparam ix42827z22479.INIT = 64'h5ACCE9163B9652AC;
    LUT6 ix42826z37260 (.O (nx42826z2), .I0 (nx42825z3), .I1 (nx42825z93), .I2 (
         nx42825z162), .I3 (nx42825z197), .I4 (nx42825z221), .I5 (nx42825z237)
         ) ;
         defparam ix42826z37260.INIT = 64'h6C5AA16DBAC58C69;
    LUT6 ix42825z39410 (.O (nx42825z2), .I0 (nx42825z3), .I1 (nx42825z93), .I2 (
         nx42825z162), .I3 (nx42825z197), .I4 (nx42825z221), .I5 (nx42825z237)
         ) ;
         defparam ix42825z39410.INIT = 64'hAE45C3B853A894CF;
    LUT6 ix42825z39995 (.O (nx42825z237), .I0 (\p_key_samp(39)  ), .I1 (
         nx42825z238), .I2 (px3060), .I3 (px2893), .I4 (px2720), .I5 (
         nx42825z242)) ;
         defparam ix42825z39995.INIT = 64'h9669699669969669;
    LUT6 ix42825z29353 (.O (nx42825z242), .I0 (nx42825z243), .I1 (px2558), .I2 (
         px2557), .I3 (px2555), .I4 (nx42825z249), .I5 (px2551)) ;
         defparam ix42825z29353.INIT = 64'h4967B59C931A6CD2;
    LUT6 ix29862z52022 (.O (px2552), .I0 (nx42825z99), .I1 (px2623), .I2 (px2622
         ), .I3 (px2621), .I4 (nx42825z119), .I5 (px2618)) ;
         defparam ix29862z52022.INIT = 64'h966352AD39D7C614;
    LUT6 ix42825z28529 (.O (nx42825z249), .I0 (\p_key_samp(35)  ), .I1 (
         nx42825z250), .I2 (nx12903z279), .I3 (nx12903z348), .I4 (nx42825z133), 
         .I5 (nx42825z251)) ;
         defparam ix42825z28529.INIT = 64'h6996966996696996;
    LUT6 ix42825z27375 (.O (nx42825z251), .I0 (nx42825z142), .I1 (nx42825z155), 
         .I2 (px2646), .I3 (px2644), .I4 (px2643), .I5 (px2642)) ;
         defparam ix42825z27375.INIT = 64'h9863C3BE69376512;
    LUT6 ix29858z47755 (.O (px2556), .I0 (px2638), .I1 (px2637), .I2 (
         nx42825z172), .I3 (px2634), .I4 (nx42825z176), .I5 (px2630)) ;
         defparam ix29858z47755.INIT = 64'hA356C9B8C235B569;
    LUT6 ix42825z28526 (.O (nx42825z243), .I0 (\p_key_samp(49)  ), .I1 (
         nx42825z244), .I2 (nx12903z277), .I3 (nx12903z336), .I4 (nx42825z129), 
         .I5 (nx42825z245)) ;
         defparam ix42825z28526.INIT = 64'h6996966996696996;
    LUT6 ix42825z59744 (.O (nx42825z245), .I0 (px2731), .I1 (px2709), .I2 (
         px2719), .I3 (nx12903z2), .I4 (nx12903z391), .I5 (px2765)) ;
         defparam ix42825z59744.INIT = 64'hE79A54291675E386;
    LUT6 ix42825z28508 (.O (nx42825z221), .I0 (\p_key_samp(7)  ), .I1 (
         nx42825z222), .I2 (px3077), .I3 (px2871), .I4 (px2710), .I5 (
         nx42825z226)) ;
         defparam ix42825z28508.INIT = 64'h6996966996696996;
    LUT6 ix42825z39685 (.O (nx42825z226), .I0 (px2570), .I1 (px2569), .I2 (
         nx42825z229), .I3 (px2566), .I4 (nx42825z233), .I5 (px2563)) ;
         defparam ix42825z39685.INIT = 64'hC92F3AC13A95953A;
    LUT6 ix42825z28517 (.O (nx42825z233), .I0 (\p_key_samp(58)  ), .I1 (
         nx42825z234), .I2 (nx12903z235), .I3 (nx12903z442), .I4 (nx42825z152), 
         .I5 (nx42825z235)) ;
         defparam ix42825z28517.INIT = 64'h6996966996696996;
    LUT6 ix42825z35102 (.O (nx42825z235), .I0 (nx12903z391), .I1 (px2709), .I2 (
         px2765), .I3 (px2719), .I4 (px2731), .I5 (nx12903z2)) ;
         defparam ix42825z35102.INIT = 64'hA6AD78D16E92834D;
    LUT6 ix42825z28514 (.O (nx42825z229), .I0 (\p_key_samp(43)  ), .I1 (
         nx42825z230), .I2 (nx12903z232), .I3 (nx12903z447), .I4 (nx42825z147), 
         .I5 (nx42825z231)) ;
         defparam ix42825z28514.INIT = 64'h6996966996696996;
    LUT6 ix42825z48017 (.O (nx42825z231), .I0 (px2621), .I1 (px2623), .I2 (
         px2622), .I3 (nx42825z119), .I4 (nx42825z99), .I5 (px2618)) ;
         defparam ix42825z48017.INIT = 64'hA739C836483EB5C3;
    LUT6 ix42825z39967 (.O (nx42825z197), .I0 (\p_key_samp(5)  ), .I1 (
         nx42825z198), .I2 (px3090), .I3 (px2881), .I4 (px2732), .I5 (
         nx42825z200)) ;
         defparam ix42825z39967.INIT = 64'h9669699669969669;
    LUT6 ix42825z24797 (.O (nx42825z200), .I0 (px2582), .I1 (nx42825z202), .I2 (
         px2579), .I3 (nx42825z206), .I4 (px2575), .I5 (px2573)) ;
         defparam ix42825z24797.INIT = 64'hDE2891CB66D65B24;
    LUT6 ix27866z29364 (.O (px2574), .I0 (nx42825z99), .I1 (px2623), .I2 (px2622
         ), .I3 (px2621), .I4 (nx42825z119), .I5 (px2618)) ;
         defparam ix27866z29364.INIT = 64'hB728847BE91C6D92;
    LUT6 ix27864z43612 (.O (px2576), .I0 (nx42825z11), .I1 (nx42825z40), .I2 (
         px2672), .I3 (px2670), .I4 (px2669), .I5 (px2668)) ;
         defparam ix27864z43612.INIT = 64'h936C96C95A96A53A;
    LUT6 ix42825z39974 (.O (nx42825z206), .I0 (\p_key_samp(12)  ), .I1 (
         nx42825z207), .I2 (nx12903z363), .I3 (nx12903z436), .I4 (nx42825z114), 
         .I5 (nx42825z208)) ;
         defparam ix42825z39974.INIT = 64'h9669699669969669;
    LUT6 ix42825z40072 (.O (nx42825z208), .I0 (nx42825z209), .I1 (px2608), .I2 (
         px2605), .I3 (px2607), .I4 (px2606), .I5 (nx42825z216)) ;
         defparam ix42825z40072.INIT = 64'h9C6372A5631E96C9;
    LUT6 ix42825z28496 (.O (nx42825z202), .I0 (\p_key_samp(21)  ), .I1 (
         nx42825z203), .I2 (nx12903z360), .I3 (nx12903z430), .I4 (nx42825z111), 
         .I5 (nx42825z204)) ;
         defparam ix42825z28496.INIT = 64'h6996966996696996;
    LUT6 ix42825z26454 (.O (nx42825z204), .I0 (nx42825z185), .I1 (px2694), .I2 (
         nx42825z189), .I3 (px2683), .I4 (px2682), .I5 (px2680)) ;
         defparam ix42825z26454.INIT = 64'h343CE666CB96619A;
    LUT6 ix42825z39944 (.O (nx42825z162), .I0 (\p_key_samp(46)  ), .I1 (
         nx42825z163), .I2 (px3136), .I3 (px2927), .I4 (px2766), .I5 (
         nx42825z166)) ;
         defparam ix42825z39944.INIT = 64'h9669699669969669;
    LUT6 ix42825z37461 (.O (nx42825z166), .I0 (nx42825z167), .I1 (px2593), .I2 (
         px2591), .I3 (nx42825z182), .I4 (px2587), .I5 (px2585)) ;
         defparam ix42825z37461.INIT = 64'hC63A29E5699D8CB2;
    LUT6 ix26867z46821 (.O (px2586), .I0 (nx42825z71), .I1 (px2654), .I2 (
         nx42825z85), .I3 (px2656), .I4 (px2658), .I5 (px2664)) ;
         defparam ix26867z46821.INIT = 64'hB4494BB86CB6B1C3;
    LUT6 ix26865z26798 (.O (px2588), .I0 (nx42825z11), .I1 (nx42825z40), .I2 (
         px2672), .I3 (px2670), .I4 (px2669), .I5 (px2668)) ;
         defparam ix26865z26798.INIT = 64'hCA2535D39C73638C;
    LUT6 ix42825z28483 (.O (nx42825z182), .I0 (\p_key_samp(52)  ), .I1 (
         nx42825z183), .I2 (nx12903z177), .I3 (nx12903z289), .I4 (nx42825z55), .I5 (
         nx42825z184)) ;
         defparam ix42825z28483.INIT = 64'h6996966996696996;
    LUT6 ix42825z27778 (.O (nx42825z184), .I0 (nx42825z185), .I1 (px2694), .I2 (
         nx42825z189), .I3 (px2683), .I4 (px2682), .I5 (px2680)) ;
         defparam ix42825z27778.INIT = 64'hE21D659A962C66D3;
    LUT6 ix25874z51339 (.O (px2592), .I0 (px2642), .I1 (px2646), .I2 (
         nx42825z142), .I3 (nx42825z155), .I4 (px2644), .I5 (px2643)) ;
         defparam ix25874z51339.INIT = 64'hDA68359A3C87C369;
    LUT6 ix25872z41477 (.O (px2594), .I0 (px2607), .I1 (px2608), .I2 (
         nx42825z209), .I3 (px2605), .I4 (nx42825z216), .I5 (px2606)) ;
         defparam ix25872z41477.INIT = 64'hD40FBA4963D09CE3;
    LUT6 ix42825z39949 (.O (nx42825z167), .I0 (\p_key_samp(10)  ), .I1 (
         nx42825z168), .I2 (nx12903z175), .I3 (nx12903z266), .I4 (nx42825z48), .I5 (
         nx42825z169)) ;
         defparam ix42825z39949.INIT = 64'h9669699669969669;
    LUT6 ix42825z40923 (.O (nx42825z169), .I0 (px2638), .I1 (px2637), .I2 (
         nx42825z172), .I3 (px2634), .I4 (nx42825z176), .I5 (px2630)) ;
         defparam ix42825z40923.INIT = 64'h69A7A31C476C9A35;
    LUT6 ix42825z28418 (.O (nx42825z93), .I0 (\p_key_samp(22)  ), .I1 (
         nx42825z94), .I2 (nx12903z344), .I3 (nx12903z393), .I4 (nx12903z414), .I5 (
         nx42825z95)) ;
         defparam ix42825z28418.INIT = 64'h6996966996696996;
    LUT6 ix42825z54175 (.O (nx42825z95), .I0 (nx42825z96), .I1 (px2615), .I2 (
         px2613), .I3 (px2611), .I4 (px2601), .I5 (nx42825z139)) ;
         defparam ix42825z54175.INIT = 64'h3EA569CAA354CE31;
    LUT6 ix42825z28452 (.O (nx42825z139), .I0 (\p_key_samp(46)  ), .I1 (
         nx42825z140), .I2 (nx12903z246), .I3 (nx12903z411), .I4 (nx12903z454), 
         .I5 (nx42825z141)) ;
         defparam ix42825z28452.INIT = 64'h6996966996696996;
    LUT6 ix42825z16214 (.O (nx42825z141), .I0 (nx42825z142), .I1 (nx42825z155), 
         .I2 (px2646), .I3 (px2644), .I4 (px2643), .I5 (px2642)) ;
         defparam ix42825z16214.INIT = 64'h3CA5D615C35A39C6;
    LUT6 ix23878z12041 (.O (px2602), .I0 (nx42825z209), .I1 (px2608), .I2 (
         px2607), .I3 (px2606), .I4 (px2605), .I5 (nx42825z216)) ;
         defparam ix23878z12041.INIT = 64'hD4E16A1C9B4C29E7;
    LUT6 ix42825z39980 (.O (nx42825z216), .I0 (\p_key_samp(60)  ), .I1 (
         nx42825z217), .I2 (nx12903z160), .I3 (nx12903z242), .I4 (nx12903z478), 
         .I5 (nx42825z218)) ;
         defparam ix42825z39980.INIT = 64'h9669699669969669;
    LUT6 ix42825z54262 (.O (nx42825z218), .I0 (px2751), .I1 (px2764), .I2 (
         nx12903z452), .I3 (nx12903z416), .I4 (nx12903z466), .I5 (nx12903z480)
         ) ;
         defparam ix42825z54262.INIT = 64'h2D2D53E8E295CE31;
    LUT6 ix42825z28502 (.O (nx42825z209), .I0 (\p_key_samp(41)  ), .I1 (
         nx42825z210), .I2 (nx12903z163), .I3 (nx12903z228), .I4 (nx12903z473), 
         .I5 (nx42825z211)) ;
         defparam ix42825z28502.INIT = 64'h6996966996696996;
    LUT6 ix42825z27502 (.O (nx42825z211), .I0 (nx42825z149), .I1 (nx42825z153), 
         .I2 (nx42825z145), .I3 (nx42825z150), .I4 (px2712), .I5 (px2711)) ;
         defparam ix42825z27502.INIT = 64'h4E939A56A69365AC;
    LUT6 ix22881z32136 (.O (px2612), .I0 (nx42825z185), .I1 (px2694), .I2 (
         nx42825z189), .I3 (px2683), .I4 (px2682), .I5 (px2680)) ;
         defparam ix22881z32136.INIT = 64'h695B872C1DB47866;
    LUT6 ix22879z51416 (.O (px2614), .I0 (px2664), .I1 (nx42825z71), .I2 (
         nx42825z85), .I3 (px2658), .I4 (px2656), .I5 (px2654)) ;
         defparam ix22879z51416.INIT = 64'hC619B1463AE9C3B6;
    LUT6 ix42825z28421 (.O (nx42825z96), .I0 (\p_key_samp(39)  ), .I1 (
         nx42825z97), .I2 (nx12903z244), .I3 (nx12903z396), .I4 (nx12903z418), .I5 (
         nx42825z98)) ;
         defparam ix42825z28421.INIT = 64'h6996966996696996;
    LUT6 ix42825z26319 (.O (nx42825z98), .I0 (nx42825z99), .I1 (px2623), .I2 (
         px2622), .I3 (px2621), .I4 (nx42825z119), .I5 (px2618)) ;
         defparam ix42825z26319.INIT = 64'h741E1EE19B61615E;
    LUT6 ix42825z28439 (.O (nx42825z119), .I0 (\p_key_samp(36)  ), .I1 (
         nx42825z120), .I2 (nx12903z145), .I3 (nx12903z405), .I4 (nx12903z422), 
         .I5 (nx42825z121)) ;
         defparam ix42825z28439.INIT = 64'h6996966996696996;
    LUT6 ix42825z55216 (.O (nx42825z121), .I0 (nx42825z122), .I1 (nx42825z123), 
         .I2 (px2729), .I3 (nx42825z127), .I4 (px2723), .I5 (nx42825z131)) ;
         defparam ix42825z55216.INIT = 64'h1CF8B64327C3D22D;
    LUT6 ix42825z28424 (.O (nx42825z99), .I0 (\p_key_samp(57)  ), .I1 (
         nx42825z100), .I2 (nx12903z147), .I3 (nx12903z401), .I4 (nx12903z426), 
         .I5 (nx42825z101)) ;
         defparam ix42825z28424.INIT = 64'h6996966996696996;
    LUT6 ix42825z6982 (.O (nx42825z101), .I0 (px2741), .I1 (nx42825z103), .I2 (
         nx42825z106), .I3 (nx42825z109), .I4 (nx42825z112), .I5 (px2733)) ;
         defparam ix42825z6982.INIT = 64'h7497E14A8B6E15D2;
    LUT6 ix42825z39821 (.O (nx42825z3), .I0 (\p_key_samp(61)  ), .I1 (nx12903z13
         ), .I2 (nx42825z4), .I3 (nx12903z126), .I4 (nx12903z211), .I5 (
         nx42825z5)) ;
         defparam ix42825z39821.INIT = 64'h9669699669969669;
    LUT6 ix42825z39151 (.O (nx42825z5), .I0 (px2706), .I1 (px2678), .I2 (
         nx42825z8), .I3 (nx42825z67), .I4 (px2640), .I5 (px2628)) ;
         defparam ix42825z39151.INIT = 64'h9BE6745A5C0393C9;
    LUT6 ix21877z43070 (.O (px2629), .I0 (px2638), .I1 (px2637), .I2 (
         nx42825z172), .I3 (px2634), .I4 (nx42825z176), .I5 (px2630)) ;
         defparam ix21877z43070.INIT = 64'hB89365CA69A7A31C;
    LUT6 ix44815z27251 (.O (px2631), .I0 (nx42825z74), .I1 (px2703), .I2 (px2702
         ), .I3 (nx42825z79), .I4 (nx42825z82), .I5 (px2698)) ;
         defparam ix44815z27251.INIT = 64'h579A98A3E93E6542;
    LUT6 ix42825z39955 (.O (nx42825z176), .I0 (\p_key_samp(5)  ), .I1 (
         nx42825z177), .I2 (nx12903z121), .I3 (nx12903z271), .I4 (nx42825z38), .I5 (
         nx42825z178)) ;
         defparam ix42825z39955.INIT = 64'h9669699669969669;
    LUT6 ix42825z22843 (.O (nx42825z178), .I0 (px2729), .I1 (nx42825z123), .I2 (
         nx42825z122), .I3 (nx42825z127), .I4 (px2723), .I5 (nx42825z131)) ;
         defparam ix42825z22843.INIT = 64'h1F61A07CAC78538F;
    LUT6 ix42825z39952 (.O (nx42825z172), .I0 (\p_key_samp(61)  ), .I1 (
         nx42825z173), .I2 (nx12903z123), .I3 (nx12903z284), .I4 (nx42825z32), .I5 (
         nx42825z174)) ;
         defparam ix42825z39952.INIT = 64'h9669699669969669;
    LUT6 ix42825z17467 (.O (nx42825z174), .I0 (px2827), .I1 (px2867), .I2 (
         nx12903z318), .I3 (nx12903z213), .I4 (px2801), .I5 (nx12903z376)) ;
         defparam ix42825z17467.INIT = 64'h6A94C56B94673E92;
    LUT6 ix43824z15348 (.O (px2639), .I0 (nx42825z14), .I1 (nx42825z17), .I2 (
         nx42825z18), .I3 (nx42825z19), .I4 (nx42825z22), .I5 (nx42825z25)) ;
         defparam ix43824z15348.INIT = 64'h61B6E92CC99636C3;
    LUT6 ix19891z57221 (.O (px2641), .I0 (nx42825z142), .I1 (nx42825z155), .I2 (
         px2646), .I3 (px2644), .I4 (px2643), .I5 (px2642)) ;
         defparam ix19891z57221.INIT = 64'h7247853CA59CDA63;
    LUT6 ix43824z45640 (.O (px2645), .I0 (nx42825z49), .I1 (nx42825z53), .I2 (
         nx42825z46), .I3 (nx42825z43), .I4 (nx42825z56), .I5 (nx42825z59)) ;
         defparam ix43824z45640.INIT = 64'h845E72C47AB1AD1B;
    LUT6 ix43820z24523 (.O (px2647), .I0 (px2764), .I1 (nx12903z416), .I2 (
         px2751), .I3 (nx12903z452), .I4 (nx12903z466), .I5 (nx12903z480)) ;
         defparam ix43820z24523.INIT = 64'h933666C96D985AA5;
    LUT6 ix42825z28466 (.O (nx42825z155), .I0 (\p_key_samp(6)  ), .I1 (
         nx42825z156), .I2 (nx12903z107), .I3 (nx12903z356), .I4 (nx12903z461), 
         .I5 (nx42825z157)) ;
         defparam ix42825z28466.INIT = 64'h6996966996696996;
    LUT6 ix42825z15868 (.O (nx42825z157), .I0 (nx42825z112), .I1 (nx42825z103), 
         .I2 (nx42825z106), .I3 (px2741), .I4 (nx42825z109), .I5 (px2733)) ;
         defparam ix42825z15868.INIT = 64'h4A7D6781876A385E;
    LUT6 ix42825z28455 (.O (nx42825z142), .I0 (\p_key_samp(7)  ), .I1 (
         nx42825z143), .I2 (nx12903z111), .I3 (nx12903z352), .I4 (nx12903z458), 
         .I5 (nx42825z144)) ;
         defparam ix42825z28455.INIT = 64'h6996966996696996;
    LUT6 ix42825z55232 (.O (nx42825z144), .I0 (nx42825z145), .I1 (px2711), .I2 (
         nx42825z149), .I3 (nx42825z150), .I4 (nx42825z153), .I5 (px2712)) ;
         defparam ix42825z55232.INIT = 64'h566A39C6A754D22D;
    LUT6 ix42825z39876 (.O (nx42825z67), .I0 (\p_key_samp(57)  ), .I1 (
         nx42825z68), .I2 (nx12903z61), .I3 (nx12903z187), .I4 (nx12903z320), .I5 (
         nx42825z69)) ;
         defparam ix42825z39876.INIT = 64'h9669699669969669;
    LUT6 ix42825z8497 (.O (nx42825z69), .I0 (px2664), .I1 (nx42825z71), .I2 (
         nx42825z85), .I3 (px2658), .I4 (px2656), .I5 (px2654)) ;
         defparam ix42825z8497.INIT = 64'hE1ADE41B66621BD4;
    LUT6 ix44815z35912 (.O (px2655), .I0 (px2729), .I1 (nx42825z123), .I2 (
         nx42825z122), .I3 (nx42825z127), .I4 (px2723), .I5 (nx42825z131)) ;
         defparam ix44815z35912.INIT = 64'h692CC2DB96F1871C;
    LUT6 ix44815z19430 (.O (px2657), .I0 (nx42825z112), .I1 (nx42825z106), .I2 (
         nx42825z103), .I3 (px2741), .I4 (nx42825z109), .I5 (px2733)) ;
         defparam ix44815z19430.INIT = 64'h346EC956DA8146BE;
    LUT6 ix44819z24282 (.O (px2659), .I0 (px2867), .I1 (nx12903z213), .I2 (
         px2827), .I3 (nx12903z318), .I4 (px2801), .I5 (nx12903z376)) ;
         defparam ix44819z24282.INIT = 64'h72A76929C29D59A6;
    LUT6 ix42825z28415 (.O (nx42825z85), .I0 (\p_key_samp(27)  ), .I1 (
         nx42825z86), .I2 (nx12903z65), .I3 (nx12903z191), .I4 (nx12903z323), .I5 (
         nx42825z87)) ;
         defparam ix42825z28415.INIT = 64'h6996966996696996;
    LUT6 ix42825z32813 (.O (nx42825z87), .I0 (nx42825z43), .I1 (nx42825z59), .I2 (
         nx42825z49), .I3 (nx42825z56), .I4 (nx42825z46), .I5 (nx42825z53)) ;
         defparam ix42825z32813.INIT = 64'h55B6A559832D7AC2;
    LUT6 ix42825z39879 (.O (nx42825z71), .I0 (\p_key_samp(42)  ), .I1 (
         nx42825z72), .I2 (nx12903z63), .I3 (nx12903z194), .I4 (nx12903z374), .I5 (
         nx42825z73)) ;
         defparam ix42825z39879.INIT = 64'h9669699669969669;
    LUT6 ix42825z33524 (.O (nx42825z73), .I0 (nx42825z74), .I1 (px2703), .I2 (
         px2702), .I3 (nx42825z79), .I4 (nx42825z82), .I5 (px2698)) ;
         defparam ix42825z33524.INIT = 64'hC52BB668825D7D94;
    LUT6 ix44819z28103 (.O (px2665), .I0 (nx42825z18), .I1 (nx42825z19), .I2 (
         nx42825z14), .I3 (nx42825z22), .I4 (nx42825z25), .I5 (nx42825z17)) ;
         defparam ix44819z28103.INIT = 64'h3CC38769DA35689A;
    LUT6 ix42825z28349 (.O (nx42825z8), .I0 (\p_key_samp(9)  ), .I1 (nx42825z9)
         , .I2 (nx12903z94), .I3 (nx12903z131), .I4 (nx12903z215), .I5 (
         nx42825z10)) ;
         defparam ix42825z28349.INIT = 64'h6996966996696996;
    LUT6 ix42825z16789 (.O (nx42825z10), .I0 (nx42825z11), .I1 (nx42825z40), .I2 (
         px2672), .I3 (px2670), .I4 (px2669), .I5 (px2668)) ;
         defparam ix42825z16789.INIT = 64'hC95AA35539A33C6C;
    LUT6 ix43816z16021 (.O (px2671), .I0 (px2867), .I1 (nx12903z213), .I2 (
         px2827), .I3 (nx12903z318), .I4 (px2801), .I5 (nx12903z376)) ;
         defparam ix43816z16021.INIT = 64'hCBA9A45987763961;
    LUT6 ix43816z59475 (.O (px2673), .I0 (nx42825z74), .I1 (px2703), .I2 (px2702
         ), .I3 (nx42825z79), .I4 (nx42825z82), .I5 (px2698)) ;
         defparam ix43816z59475.INIT = 64'h61163DDA61CBE31C;
    LUT6 ix42825z28378 (.O (nx42825z40), .I0 (\p_key_samp(23)  ), .I1 (
         nx42825z41), .I2 (nx12903z101), .I3 (nx12903z171), .I4 (nx12903z262), .I5 (
         nx42825z42)) ;
         defparam ix42825z28378.INIT = 64'h6996966996696996;
    LUT6 ix42825z9240 (.O (nx42825z42), .I0 (nx42825z43), .I1 (nx42825z46), .I2 (
         nx42825z49), .I3 (nx42825z53), .I4 (nx42825z56), .I5 (nx42825z59)) ;
         defparam ix42825z9240.INIT = 64'h3E61E11E61971ED2;
    LUT6 ix42825z28352 (.O (nx42825z11), .I0 (\p_key_samp(30)  ), .I1 (
         nx42825z12), .I2 (nx12903z99), .I3 (nx12903z135), .I4 (nx12903z305), .I5 (
         nx42825z13)) ;
         defparam ix42825z28352.INIT = 64'h6996966996696996;
    LUT6 ix42825z41937 (.O (nx42825z13), .I0 (nx42825z14), .I1 (nx42825z17), .I2 (
         nx42825z18), .I3 (nx42825z19), .I4 (nx42825z22), .I5 (nx42825z25)) ;
         defparam ix42825z41937.INIT = 64'h3C87D2A983789EA5;
    LUT6 ix16892z12698 (.O (px2679), .I0 (nx42825z185), .I1 (px2694), .I2 (
         nx42825z189), .I3 (px2683), .I4 (px2682), .I5 (px2680)) ;
         defparam ix16892z12698.INIT = 64'hAC69D187731D2C78;
    LUT6 ix45810z16839 (.O (px2681), .I0 (px2764), .I1 (nx12903z416), .I2 (
         px2751), .I3 (nx12903z452), .I4 (nx12903z466), .I5 (nx12903z480)) ;
         defparam ix45810z16839.INIT = 64'h865E782DC3E13C96;
    LUT6 ix42825z28489 (.O (nx42825z189), .I0 (\p_key_samp(19)  ), .I1 (
         nx42825z190), .I2 (nx12903z51), .I3 (nx12903z300), .I4 (nx12903z389), .I5 (
         nx42825z191)) ;
         defparam ix42825z28489.INIT = 64'h6996966996696996;
    LUT6 ix42825z60784 (.O (nx42825z191), .I0 (nx42825z14), .I1 (nx42825z17), .I2 (
         nx42825z18), .I3 (nx42825z19), .I4 (nx42825z22), .I5 (nx42825z25)) ;
         defparam ix42825z60784.INIT = 64'hE52690C11AC5E7BB;
    LUT6 ix42825z39841 (.O (nx42825z25), .I0 (\p_key_samp(55)  ), .I1 (
         nx42825z26), .I2 (nx12903z58), .I3 (nx12903z139), .I4 (nx12903z311), .I5 (
         nx42825z27)) ;
         defparam ix42825z39841.INIT = 64'h9669699669969669;
    LUT6 ix42825z37836 (.O (nx42825z27), .I0 (px2812), .I1 (px2810), .I2 (
         nx42825z30), .I3 (nx42825z33), .I4 (nx42825z36), .I5 (px2803)) ;
         defparam ix42825z37836.INIT = 64'hDA61718DB5478E92;
    LUT6 ix42825z28363 (.O (nx42825z22), .I0 (\p_key_samp(37)  ), .I1 (px3322), 
         .I2 (px3321), .I3 (px3095), .I4 (px2885), .I5 (px2734)) ;
         defparam ix42825z28363.INIT = 64'h6996966996696996;
    LUT6 ix42825z28360 (.O (nx42825z19), .I0 (\p_key_samp(23)  ), .I1 (px3316), 
         .I2 (px3315), .I3 (px3092), .I4 (px2891), .I5 (px2742)) ;
         defparam ix42825z28360.INIT = 64'h6996966996696996;
    LUT6 ix42825z28359 (.O (nx42825z18), .I0 (\p_key_samp(46)  ), .I1 (px3723), 
         .I2 (px3504), .I3 (px3281), .I4 (px3058), .I5 (px2869)) ;
         defparam ix42825z28359.INIT = 64'h6996966996696996;
    LUT6 ix42825z39833 (.O (nx42825z17), .I0 (\p_key_samp(13)  ), .I1 (
         nx12903z467), .I2 (px3359), .I3 (px3119), .I4 (px2914), .I5 (px2748)) ;
         defparam ix42825z39833.INIT = 64'h9669699669969669;
    LUT6 ix42825z28355 (.O (nx42825z14), .I0 (\p_key_samp(20)  ), .I1 (
         nx42825z15), .I2 (nx12903z55), .I3 (nx12903z137), .I4 (nx12903z308), .I5 (
         nx42825z16)) ;
         defparam ix42825z28355.INIT = 64'h6996966996696996;
    LUT6 ix42825z15812 (.O (nx42825z16), .I0 (nx12903z321), .I1 (px2823), .I2 (
         px2821), .I3 (nx12903z326), .I4 (nx12903z330), .I5 (nx12903z372)) ;
         defparam ix42825z15812.INIT = 64'h689DC75A97A13895;
    LUT6 ix45810z39347 (.O (px2695), .I0 (nx42825z150), .I1 (nx42825z149), .I2 (
         nx42825z145), .I3 (px2711), .I4 (px2712), .I5 (nx42825z153)) ;
         defparam ix45810z39347.INIT = 64'hC61B6B3C4BB4948B;
    LUT6 ix42825z28486 (.O (nx42825z185), .I0 (\p_key_samp(33)  ), .I1 (
         nx42825z186), .I2 (nx12903z27), .I3 (nx12903z294), .I4 (nx12903z382), .I5 (
         nx42825z187)) ;
         defparam ix42825z28486.INIT = 64'h6996966996696996;
    LUT6 ix42825z57623 (.O (nx42825z187), .I0 (nx42825z74), .I1 (px2703), .I2 (
         px2702), .I3 (nx42825z79), .I4 (nx42825z82), .I5 (px2698)) ;
         defparam ix42825z57623.INIT = 64'hD34921BE2856DB65;
    LUT6 ix42825z28413 (.O (nx42825z82), .I0 (\p_key_samp(47)  ), .I1 (
         nx12903z252), .I2 (nx32966z9), .I3 (nx12903z196), .I4 (nx12903z253), .I5 (
         nx42825z83)) ;
         defparam ix42825z28413.INIT = 64'h6996966996696996;
    LUT6 ix42825z17090 (.O (nx42825z83), .I0 (nx12903z260), .I1 (nx12903z217), .I2 (
         px2866), .I3 (px2841), .I4 (nx12903z257), .I5 (nx12903z303)) ;
         defparam ix42825z17090.INIT = 64'hCD3253A896C53D5A;
    LUT6 ix42825z39885 (.O (nx42825z79), .I0 (\p_key_samp(30)  ), .I1 (px3305), 
         .I2 (px3304), .I3 (px3068), .I4 (px2899), .I5 (px2730)) ;
         defparam ix42825z39885.INIT = 64'h9669699669969669;
    LUT6 ix42825z39882 (.O (nx42825z74), .I0 (\p_key_samp(21)  ), .I1 (
         nx42825z75), .I2 (nx32966z7), .I3 (nx12903z200), .I4 (nx12903z224), .I5 (
         nx42825z76)) ;
         defparam ix42825z39882.INIT = 64'h9669699669969669;
    LUT6 ix42825z56278 (.O (nx42825z76), .I0 (px2780), .I1 (nx12903z471), .I2 (
         px2777), .I3 (nx12903z475), .I4 (nx12903z476), .I5 (px2773)) ;
         defparam ix42825z56278.INIT = 64'h66E9A590922DD673;
    LUT6 ix12904z50833 (.O (px2707), .I0 (nx12903z391), .I1 (px2765), .I2 (
         px2719), .I3 (px2731), .I4 (px2709), .I5 (nx12903z2)) ;
         defparam ix12904z50833.INIT = 64'hD9843D526635C16F;
    LUT6 ix12903z61247 (.O (px2708), .I0 (nx12903z2), .I1 (px2765), .I2 (
         nx12903z391), .I3 (px2731), .I4 (px2719), .I5 (px2709)) ;
         defparam ix12903z61247.INIT = 64'hCA3C30D675A2EA1D;
    LUT6 ix42825z52991 (.O (px2710), .I0 (nx42825z149), .I1 (nx42825z153), .I2 (
         nx42825z145), .I3 (nx42825z150), .I4 (px2712), .I5 (px2711)) ;
         defparam ix42825z52991.INIT = 64'h9A3507DA35C9C935;
    LUT6 ix42825z39937 (.O (nx42825z150), .I0 (\p_key_samp(26)  ), .I1 (
         nx42825z151), .I2 (nx12903z20), .I3 (nx12903z235), .I4 (nx12903z442), .I5 (
         nx42825z152)) ;
         defparam ix42825z39937.INIT = 64'h9669699669969669;
    LUT6 ix42825z36989 (.O (nx42825z152), .I0 (nx61487z5), .I1 (px2926), .I2 (
         nx61487z2), .I3 (px2870), .I4 (px2892), .I5 (nx61487z8)) ;
         defparam ix42825z36989.INIT = 64'h55E9691DC3168AE3;
    LUT6 ix42825z28458 (.O (nx42825z145), .I0 (\p_key_samp(11)  ), .I1 (
         nx42825z146), .I2 (nx12903z22), .I3 (nx12903z232), .I4 (nx12903z447), .I5 (
         nx42825z147)) ;
         defparam ix42825z28458.INIT = 64'h6996966996696996;
    LUT6 ix42825z9335 (.O (nx42825z147), .I0 (px2760), .I1 (nx12903z420), .I2 (
         nx12903z437), .I3 (nx12903z424), .I4 (px2763), .I5 (nx12903z450)) ;
         defparam ix42825z9335.INIT = 64'hE7C82936C83D1EE1;
    LUT6 ix42825z39940 (.O (nx42825z153), .I0 (\p_key_samp(60)  ), .I1 (
         nx42825z50), .I2 (px3338), .I3 (px3160), .I4 (px2945), .I5 (px2786)) ;
         defparam ix42825z39940.INIT = 64'h9669699669969669;
    LUT6 ix42825z39936 (.O (nx42825z149), .I0 (\p_key_samp(49)  ), .I1 (
         nx12903z377), .I2 (px3408), .I3 (px3245), .I4 (px2985), .I5 (px2790)) ;
         defparam ix42825z39936.INIT = 64'h9669699669969669;
    LUT6 ix42825z21503 (.O (px2720), .I0 (px2729), .I1 (nx42825z123), .I2 (
         nx42825z122), .I3 (nx42825z127), .I4 (px2723), .I5 (nx42825z131)) ;
         defparam ix42825z21503.INIT = 64'h8358D4B63CE74E29;
    LUT6 ix42825z39924 (.O (nx42825z131), .I0 (\p_key_samp(3)  ), .I1 (
         nx42825z132), .I2 (nx12903z77), .I3 (nx12903z279), .I4 (nx12903z348), .I5 (
         nx42825z133)) ;
         defparam ix42825z39924.INIT = 64'h9669699669969669;
    LUT6 ix42825z13119 (.O (nx42825z133), .I0 (nx12903z463), .I1 (nx12903z455), 
         .I2 (nx12903z459), .I3 (nx12903z464), .I4 (nx12903z456), .I5 (px2835)
         ) ;
         defparam ix42825z13119.INIT = 64'h7470D26C5AC72DB2;
    LUT6 ix42825z28446 (.O (nx42825z127), .I0 (\p_key_samp(17)  ), .I1 (
         nx42825z128), .I2 (nx12903z79), .I3 (nx12903z277), .I4 (nx12903z336), .I5 (
         nx42825z129)) ;
         defparam ix42825z28446.INIT = 64'h6996966996696996;
    LUT6 ix42825z24359 (.O (nx42825z129), .I0 (nx61487z2), .I1 (px2926), .I2 (
         nx61487z5), .I3 (px2892), .I4 (nx61487z8), .I5 (px2870)) ;
         defparam ix42825z24359.INIT = 64'h69C71E69C322599D;
    LUT6 ix42825z39917 (.O (nx42825z122), .I0 (\p_key_samp(34)  ), .I1 (
         nx42825z60), .I2 (px3335), .I3 (px3151), .I4 (px2941), .I5 (px2768)) ;
         defparam ix42825z39917.INIT = 64'h9669699669969669;
    LUT6 ix42825z28443 (.O (nx42825z123), .I0 (\p_key_samp(59)  ), .I1 (px3308)
         , .I2 (px3307), .I3 (px3073), .I4 (px2895), .I5 (px2728)) ;
         defparam ix42825z28443.INIT = 64'h6996966996696996;
    LUT6 ix42825z29471 (.O (px2728), .I0 (px2763), .I1 (nx12903z420), .I2 (
         px2760), .I3 (nx12903z424), .I4 (nx12903z437), .I5 (nx12903z450)) ;
         defparam ix42825z29471.INIT = 64'hE11E59E19E946D98;
    LUT6 ix42825z60682 (.O (px2730), .I0 (px2812), .I1 (px2810), .I2 (nx42825z30
         ), .I3 (nx42825z33), .I4 (nx42825z36), .I5 (px2803)) ;
         defparam ix42825z60682.INIT = 64'hB65818EB29D1E7A4;
    LUT6 ix42825z56277 (.O (px2732), .I0 (px2741), .I1 (nx42825z103), .I2 (
         nx42825z106), .I3 (nx42825z109), .I4 (nx42825z112), .I5 (px2733)) ;
         defparam ix42825z56277.INIT = 64'h8754B9E2A14BD61D;
    LUT6 ix42825z24344 (.O (px2734), .I0 (px2763), .I1 (nx12903z420), .I2 (
         px2760), .I3 (nx12903z424), .I4 (nx12903z437), .I5 (nx12903z450)) ;
         defparam ix42825z24344.INIT = 64'h7A2C2D78B45A59E1;
    LUT6 ix42825z39911 (.O (nx42825z112), .I0 (\p_key_samp(45)  ), .I1 (
         nx42825z113), .I2 (nx12903z36), .I3 (nx12903z363), .I4 (nx12903z436), .I5 (
         nx42825z114)) ;
         defparam ix42825z39911.INIT = 64'h9669699669969669;
    LUT6 ix42825z39881 (.O (nx42825z114), .I0 (nx12903z471), .I1 (nx12903z476), 
         .I2 (px2780), .I3 (px2777), .I4 (px2773), .I5 (nx12903z475)) ;
         defparam ix42825z39881.INIT = 64'h93582DE67CA39649;
    LUT6 ix42825z39908 (.O (nx42825z109), .I0 (\p_key_samp(54)  ), .I1 (
         nx42825z110), .I2 (nx12903z31), .I3 (nx12903z360), .I4 (nx12903z430), .I5 (
         nx42825z111)) ;
         defparam ix42825z39908.INIT = 64'h9669699669969669;
    LUT6 ix42825z37366 (.O (nx42825z111), .I0 (nx12903z380), .I1 (px2797), .I2 (
         px2796), .I3 (px2794), .I4 (px2793), .I5 (nx12903z387)) ;
         defparam ix42825z37366.INIT = 64'hD99633C699258C79;
    LUT6 ix42825z39905 (.O (nx42825z106), .I0 (\p_key_samp(63)  ), .I1 (px3403)
         , .I2 (px3392), .I3 (px3187), .I4 (px2953), .I5 (px2828)) ;
         defparam ix42825z39905.INIT = 64'h9669699669969669;
    LUT6 ix42825z39902 (.O (nx42825z103), .I0 (\p_key_samp(4)  ), .I1 (px3406), 
         .I2 (px3405), .I3 (px3221), .I4 (px3057), .I5 (px2868)) ;
         defparam ix42825z39902.INIT = 64'h9669699669969669;
    LUT6 ix42825z52042 (.O (px2742), .I0 (px2866), .I1 (nx12903z217), .I2 (
         nx12903z257), .I3 (nx12903z260), .I4 (nx12903z303), .I5 (px2841)) ;
         defparam ix42825z52042.INIT = 64'h43BC2DD2B969C616;
    LUT6 ix12903z28687 (.O (nx12903z391), .I0 (\p_key_samp(63)  ), .I1 (
         nx12903z392), .I2 (nx12903z88), .I3 (nx12903z344), .I4 (nx12903z393), .I5 (
         nx12903z414)) ;
         defparam ix12903z28687.INIT = 64'h6996966996696996;
    LUT6 ix12903z37710 (.O (nx12903z414), .I0 (px2764), .I1 (nx12903z416), .I2 (
         px2751), .I3 (nx12903z452), .I4 (nx12903z466), .I5 (nx12903z480)) ;
         defparam ix12903z37710.INIT = 64'hBA6953B5453A8CC3;
    LUT6 ix12903z28759 (.O (nx12903z480), .I0 (\p_key_samp(53)  ), .I1 (px3354)
         , .I2 (px3353), .I3 (px3109), .I4 (px2907), .I5 (px2746)) ;
         defparam ix12903z28759.INIT = 64'h6996966996696996;
    LUT6 ix12903z28331 (.O (px2746), .I0 (nx12903z380), .I1 (px2797), .I2 (
         px2796), .I3 (px2794), .I4 (px2793), .I5 (nx12903z387)) ;
         defparam ix12903z28331.INIT = 64'h41B99A27BC4967E8;
    LUT6 ix12903z40223 (.O (nx12903z466), .I0 (\p_key_samp(62)  ), .I1 (
         nx12903z467), .I2 (px3359), .I3 (px3119), .I4 (px2914), .I5 (px2748)) ;
         defparam ix12903z40223.INIT = 64'h9669699669969669;
    LUT6 ix12903z20399 (.O (px2748), .I0 (px2780), .I1 (nx12903z471), .I2 (
         px2777), .I3 (nx12903z475), .I4 (nx12903z476), .I5 (px2773)) ;
         defparam ix12903z20399.INIT = 64'h9EA3B149B59448F6;
    LUT6 ix12903z40209 (.O (nx12903z452), .I0 (\p_key_samp(14)  ), .I1 (
         nx12903z453), .I2 (nx12903z46), .I3 (nx12903z246), .I4 (nx12903z411), .I5 (
         nx12903z454)) ;
         defparam ix12903z40209.INIT = 64'h9669699669969669;
    LUT6 ix12903z39459 (.O (nx12903z454), .I0 (nx12903z455), .I1 (nx12903z456), 
         .I2 (nx12903z459), .I3 (px2835), .I4 (nx12903z463), .I5 (nx12903z464)
         ) ;
         defparam ix12903z39459.INIT = 64'hB9584EA5CC879378;
    LUT6 ix7924z12005 (.O (px2752), .I0 (nx12903z321), .I1 (px2823), .I2 (px2821
         ), .I3 (nx12903z326), .I4 (nx12903z330), .I5 (nx12903z372)) ;
         defparam ix7924z12005.INIT = 64'hE549913C7E9629C3;
    LUT6 ix12903z28706 (.O (nx12903z416), .I0 (\p_key_samp(7)  ), .I1 (
         nx12903z417), .I2 (nx12903z41), .I3 (nx12903z244), .I4 (nx12903z396), .I5 (
         nx12903z418)) ;
         defparam ix12903z28706.INIT = 64'h6996966996696996;
    LUT6 ix12903z17204 (.O (nx12903z418), .I0 (px2763), .I1 (nx12903z420), .I2 (
         px2760), .I3 (nx12903z424), .I4 (nx12903z437), .I5 (nx12903z450)) ;
         defparam ix12903z17204.INIT = 64'h2CB6C359926D3CA6;
    LUT6 ix12903z40208 (.O (nx12903z450), .I0 (\p_key_samp(2)  ), .I1 (
         nx12903z327), .I2 (px3460), .I3 (px3232), .I4 (px2973), .I5 (px2820)) ;
         defparam ix12903z40208.INIT = 64'h9669699669969669;
    LUT6 ix12903z28722 (.O (nx12903z437), .I0 (\p_key_samp(11)  ), .I1 (px3422)
         , .I2 (px3421), .I3 (px3278), .I4 (px2997), .I5 (px2798)) ;
         defparam ix12903z28722.INIT = 64'h6996966996696996;
    LUT6 ix12903z28712 (.O (nx12903z424), .I0 (\p_key_samp(25)  ), .I1 (
         nx12903z425), .I2 (nx337z6), .I3 (nx12903z147), .I4 (nx12903z401), .I5 (
         nx12903z426)) ;
         defparam ix12903z28712.INIT = 64'h6996966996696996;
    LUT6 ix12903z26913 (.O (nx12903z426), .I0 (px2890), .I1 (nx12903z428), .I2 (
         px2887), .I3 (px2886), .I4 (px2884), .I5 (nx12903z434)) ;
         defparam ix12903z26913.INIT = 64'hEB2935D66453628D;
    LUT6 ix45810z28353 (.O (nx45810z10), .I0 (\plaintext(8)  ), .I1 (nx34235z25)
         , .I2 (nx24265z31), .I3 (nx337z6), .I4 (nx12903z147), .I5 (nx12903z401)
         ) ;
         defparam ix45810z28353.INIT = 64'h6996966996696996;
    LUT6 ix12903z28709 (.O (nx12903z420), .I0 (\p_key_samp(35)  ), .I1 (
         nx12903z421), .I2 (nx337z4), .I3 (nx12903z145), .I4 (nx12903z405), .I5 (
         nx12903z422)) ;
         defparam ix12903z28709.INIT = 64'h6996966996696996;
    LUT6 ix12903z24826 (.O (nx12903z422), .I0 (nx12903z334), .I1 (nx12903z346), 
         .I2 (px2898), .I3 (px2897), .I4 (px2896), .I5 (px2894)) ;
         defparam ix12903z24826.INIT = 64'h6C923CA553AD5A69;
    LUT6 ix42825z12148 (.O (px2766), .I0 (nx42825z49), .I1 (nx42825z53), .I2 (
         nx42825z46), .I3 (nx42825z43), .I4 (nx42825z56), .I5 (nx42825z59)) ;
         defparam ix42825z12148.INIT = 64'h635A4E379C2729D2;
    LUT6 ix42825z39872 (.O (nx42825z59), .I0 (\p_key_samp(1)  ), .I1 (nx42825z60
         ), .I2 (px3335), .I3 (px3151), .I4 (px2941), .I5 (px2768)) ;
         defparam ix42825z39872.INIT = 64'h9669699669969669;
    LUT6 ix42825z44784 (.O (px2768), .I0 (px2866), .I1 (nx12903z217), .I2 (
         nx12903z257), .I3 (nx12903z260), .I4 (nx12903z303), .I5 (px2841)) ;
         defparam ix42825z44784.INIT = 64'h967A4569A55AA996;
    LUT6 ix42825z28394 (.O (nx42825z56), .I0 (\p_key_samp(27)  ), .I1 (px3333), 
         .I2 (px3332), .I3 (px3154), .I4 (px2943), .I5 (px2770)) ;
         defparam ix42825z28394.INIT = 64'h6996966996696996;
    LUT6 ix42825z16116 (.O (px2770), .I0 (nx12903z372), .I1 (nx12903z330), .I2 (
         px2821), .I3 (nx12903z321), .I4 (nx12903z326), .I5 (px2823)) ;
         defparam ix42825z16116.INIT = 64'hE21E4CE316E1399E;
    LUT6 ix42825z39856 (.O (nx42825z43), .I0 (\p_key_samp(58)  ), .I1 (px3342), 
         .I2 (px3341), .I3 (px3138), .I4 (px2929), .I5 (px2772)) ;
         defparam ix42825z39856.INIT = 64'h9669699669969669;
    LUT6 ix42825z35886 (.O (px2772), .I0 (px2780), .I1 (nx12903z471), .I2 (
         px2777), .I3 (nx12903z475), .I4 (nx12903z476), .I5 (px2773)) ;
         defparam ix42825z35886.INIT = 64'hC395999B7C0A86E5;
    LUT6 ix12903z40231 (.O (nx12903z476), .I0 (\p_key_samp(59)  ), .I1 (
         nx12903z477), .I2 (nx4319z3), .I3 (nx12903z160), .I4 (nx12903z242), .I5 (
         nx12903z478)) ;
         defparam ix12903z40231.INIT = 64'h9669699669969669;
    LUT6 ix12903z16780 (.O (nx12903z478), .I0 (nx12903z409), .I1 (nx12903z394), 
         .I2 (px2913), .I3 (px2906), .I4 (px2908), .I5 (px2912)) ;
         defparam ix12903z16780.INIT = 64'hCA355A3965633ACC;
    LUT6 ix12903z28755 (.O (nx12903z475), .I0 (\p_key_samp(27)  ), .I1 (
         nx12903z331), .I2 (px3448), .I3 (px3229), .I4 (px2970), .I5 (px2818)) ;
         defparam ix12903z28755.INIT = 64'h6996966996696996;
    LUT6 ix12903z28752 (.O (nx12903z471), .I0 (\p_key_samp(9)  ), .I1 (
         nx12903z472), .I2 (nx4319z5), .I3 (nx12903z163), .I4 (nx12903z228), .I5 (
         nx12903z473)) ;
         defparam ix12903z28752.INIT = 64'h6996966996696996;
    LUT6 ix12903z16415 (.O (nx12903z473), .I0 (px2879), .I1 (px2878), .I2 (
         px2877), .I3 (nx12903z440), .I4 (nx12903z445), .I5 (px2872)) ;
         defparam ix12903z16415.INIT = 64'hB359866C9C5A3963;
    LUT6 ix42825z39859 (.O (nx42825z46), .I0 (\p_key_samp(41)  ), .I1 (
         nx42825z47), .I2 (nx35956z4), .I3 (nx12903z175), .I4 (nx12903z266), .I5 (
         nx42825z48)) ;
         defparam ix42825z39859.INIT = 64'h9669699669969669;
    LUT6 ix42825z10986 (.O (nx42825z48), .I0 (px2812), .I1 (px2810), .I2 (
         nx42825z30), .I3 (nx42825z33), .I4 (nx42825z36), .I5 (px2803)) ;
         defparam ix42825z10986.INIT = 64'h1ADB4768EB24259E;
    LUT6 ix42825z39866 (.O (nx42825z53), .I0 (\p_key_samp(51)  ), .I1 (
         nx42825z54), .I2 (nx35956z6), .I3 (nx12903z177), .I4 (nx12903z289), .I5 (
         nx42825z55)) ;
         defparam ix42825z39866.INIT = 64'h9669699669969669;
    LUT6 ix42825z9199 (.O (nx42825z55), .I0 (nx12903z380), .I1 (px2797), .I2 (
         px2796), .I3 (px2794), .I4 (px2793), .I5 (nx12903z387)) ;
         defparam ix42825z9199.INIT = 64'h969ED261A5931E9C;
    LUT6 ix42825z39862 (.O (nx42825z49), .I0 (\p_key_samp(18)  ), .I1 (
         nx42825z50), .I2 (px3338), .I3 (px3160), .I4 (px2945), .I5 (px2786)) ;
         defparam ix42825z39862.INIT = 64'h9669699669969669;
    LUT6 ix42825z55544 (.O (px2786), .I0 (nx12903z463), .I1 (nx12903z459), .I2 (
         nx12903z464), .I3 (nx12903z455), .I4 (px2835), .I5 (nx12903z456)) ;
         defparam ix42825z55544.INIT = 64'hD22D2CD62D66D3A8;
    LUT6 ix12903z39820 (.O (nx12903z2), .I0 (\p_key_samp(37)  ), .I1 (nx12903z3)
         , .I2 (nx12903z4), .I3 (nx12903z13), .I4 (nx12903z126), .I5 (
         nx12903z211)) ;
         defparam ix12903z39820.INIT = 64'h9669699669969669;
    LUT6 ix12903z13726 (.O (nx12903z211), .I0 (px2867), .I1 (nx12903z213), .I2 (
         px2827), .I3 (nx12903z318), .I4 (px2801), .I5 (nx12903z376)) ;
         defparam ix12903z13726.INIT = 64'h6A34DC47615A2FB4;
    LUT6 ix12903z40151 (.O (nx12903z376), .I0 (\p_key_samp(43)  ), .I1 (
         nx12903z377), .I2 (px3408), .I3 (px3245), .I4 (px2985), .I5 (px2790)) ;
         defparam ix12903z40151.INIT = 64'h9669699669969669;
    LUT6 ix12903z52400 (.O (px2790), .I0 (nx12903z380), .I1 (px2797), .I2 (
         px2796), .I3 (px2794), .I4 (px2793), .I5 (nx12903z387)) ;
         defparam ix12903z52400.INIT = 64'hE41B59B22BC4C63E;
    LUT6 ix12903z28684 (.O (nx12903z387), .I0 (\p_key_samp(50)  ), .I1 (
         nx12903z388), .I2 (nx5318z9), .I3 (nx12903z51), .I4 (nx12903z300), .I5 (
         nx12903z389)) ;
         defparam ix12903z28684.INIT = 64'h6996966996696996;
    LUT6 ix12903z20237 (.O (nx12903z389), .I0 (nx12903z306), .I1 (nx12903z309), 
         .I2 (px2847), .I3 (px2846), .I4 (px2845), .I5 (px2844)) ;
         defparam ix12903z20237.INIT = 64'h9C62EB3CCD964895;
    LUT6 ix45810z35734 (.O (px2795), .I0 (nx12903z394), .I1 (px2913), .I2 (
         px2912), .I3 (nx12903z409), .I4 (px2908), .I5 (px2906)) ;
         defparam ix45810z35734.INIT = 64'h839C7D6179998666;
    LUT6 ix12903z40200 (.O (px2798), .I0 (nx12903z440), .I1 (px2877), .I2 (
         px2872), .I3 (nx12903z445), .I4 (px2878), .I5 (px2879)) ;
         defparam ix12903z40200.INIT = 64'hBC276BD0C31C966A;
    LUT6 ix12903z28681 (.O (nx12903z380), .I0 (\p_key_samp(1)  ), .I1 (
         nx12903z381), .I2 (nx5318z6), .I3 (nx12903z27), .I4 (nx12903z294), .I5 (
         nx12903z382)) ;
         defparam ix12903z28681.INIT = 64'h6996966996696996;
    LUT6 ix12903z59899 (.O (nx12903z382), .I0 (px2860), .I1 (px2858), .I2 (
         px2859), .I3 (nx12903z222), .I4 (nx12903z251), .I5 (px2865)) ;
         defparam ix12903z59899.INIT = 64'hE79A54291675E386;
    LUT6 ix1940z20169 (.O (px2802), .I0 (px2812), .I1 (px2810), .I2 (nx42825z30)
         , .I3 (nx42825z33), .I4 (nx42825z36), .I5 (px2803)) ;
         defparam ix1940z20169.INIT = 64'h86B2D15E724D49A7;
    LUT6 ix42825z39850 (.O (nx42825z36), .I0 (\p_key_samp(38)  ), .I1 (
         nx42825z37), .I2 (nx13298z60), .I3 (nx12903z121), .I4 (nx12903z271), .I5 (
         nx42825z38)) ;
         defparam ix42825z39850.INIT = 64'h9669699669969669;
    LUT6 ix42825z31469 (.O (nx42825z38), .I0 (nx12903z334), .I1 (nx12903z346), .I2 (
         px2898), .I3 (px2897), .I4 (px2896), .I5 (px2894)) ;
         defparam ix42825z31469.INIT = 64'hB6C94C331A6975AA;
    LUT6 ix42825z28372 (.O (nx42825z33), .I0 (\p_key_samp(47)  ), .I1 (px3440), 
         .I2 (px3439), .I3 (px3172), .I4 (px3022), .I5 (px2807)) ;
         defparam ix42825z28372.INIT = 64'h6996966996696996;
    LUT6 ix42825z26821 (.O (px2807), .I0 (nx12903z306), .I1 (nx12903z309), .I2 (
         px2847), .I3 (px2846), .I4 (px2845), .I5 (px2844)) ;
         defparam ix42825z26821.INIT = 64'hE2273CDA9C5A6385;
    LUT6 ix42825z28369 (.O (nx42825z30), .I0 (\p_key_samp(29)  ), .I1 (
         nx42825z31), .I2 (nx13298z70), .I3 (nx12903z123), .I4 (nx12903z284), .I5 (
         nx42825z32)) ;
         defparam ix42825z28369.INIT = 64'h6996966996696996;
    LUT6 ix42825z52827 (.O (nx42825z32), .I0 (nx12903z185), .I1 (px3056), .I2 (
         px3016), .I3 (px2984), .I4 (px2952), .I5 (nx12903z129)) ;
         defparam ix42825z52827.INIT = 64'h661B1EE1B469C91E;
    LUT6 ix44815z50847 (.O (px2811), .I0 (nx12903z251), .I1 (px2865), .I2 (
         px2859), .I3 (px2860), .I4 (nx12903z222), .I5 (px2858)) ;
         defparam ix44815z50847.INIT = 64'hD98466353D52C16F;
    LUT6 ix12903z40103 (.O (nx12903z318), .I0 (\p_key_samp(25)  ), .I1 (
         nx12903z319), .I2 (nx12903z8), .I3 (nx12903z61), .I4 (nx12903z187), .I5 (
         nx12903z320)) ;
         defparam ix12903z40103.INIT = 64'h9669699669969669;
    LUT6 ix12903z24556 (.O (nx12903z320), .I0 (nx12903z321), .I1 (px2823), .I2 (
         px2821), .I3 (nx12903z326), .I4 (nx12903z330), .I5 (nx12903z372)) ;
         defparam ix12903z24556.INIT = 64'h067CD993F20759AC;
    LUT6 ix12903z28672 (.O (nx12903z372), .I0 (\p_key_samp(10)  ), .I1 (
         nx12903z373), .I2 (nx7312z7), .I3 (nx12903z63), .I4 (nx12903z194), .I5 (
         nx12903z374)) ;
         defparam ix12903z28672.INIT = 64'h6996966996696996;
    LUT6 ix12903z40390 (.O (nx12903z374), .I0 (px2865), .I1 (nx12903z222), .I2 (
         nx12903z251), .I3 (px2860), .I4 (px2859), .I5 (px2858)) ;
         defparam ix12903z40390.INIT = 64'h9768E49BF099960D;
    LUT6 ix12903z28638 (.O (nx12903z330), .I0 (\p_key_samp(33)  ), .I1 (
         nx12903z331), .I2 (px3448), .I3 (px3229), .I4 (px2970), .I5 (px2818)) ;
         defparam ix12903z28638.INIT = 64'h6996966996696996;
    LUT6 ix12903z15527 (.O (px2818), .I0 (nx12903z334), .I1 (nx12903z346), .I2 (
         px2898), .I3 (px2897), .I4 (px2896), .I5 (px2894)) ;
         defparam ix12903z15527.INIT = 64'h1CF5E926C923365C;
    LUT6 ix12903z40109 (.O (nx12903z326), .I0 (\p_key_samp(44)  ), .I1 (
         nx12903z327), .I2 (px3460), .I3 (px3232), .I4 (px2973), .I5 (px2820)) ;
         defparam ix12903z40109.INIT = 64'h9669699669969669;
    LUT6 ix12903z35267 (.O (px2820), .I0 (px2844), .I1 (nx12903z309), .I2 (
         px2847), .I3 (nx12903z306), .I4 (px2845), .I5 (px2846)) ;
         defparam ix12903z35267.INIT = 64'h8799788779A2837C;
    LUT6 ix44815z12030 (.O (px2822), .I0 (px2890), .I1 (nx12903z428), .I2 (
         px2887), .I3 (px2886), .I4 (px2884), .I5 (nx12903z434)) ;
         defparam ix44815z12030.INIT = 64'hB19D5C62493A29D7;
    LUT6 ix44819z35752 (.O (px2824), .I0 (px2984), .I1 (px3016), .I2 (
         nx12903z185), .I3 (px3056), .I4 (px2952), .I5 (nx12903z129)) ;
         defparam ix44819z35752.INIT = 64'hE0930FE8D36C8675;
    LUT6 ix12903z28631 (.O (nx12903z321), .I0 (\p_key_samp(58)  ), .I1 (
         nx12903z322), .I2 (nx7312z3), .I3 (nx12903z65), .I4 (nx12903z191), .I5 (
         nx12903z323)) ;
         defparam ix12903z28631.INIT = 64'h6996966996696996;
    LUT6 ix12903z17413 (.O (nx12903z323), .I0 (px2940), .I1 (px2942), .I2 (
         px2944), .I3 (px2928), .I4 (nx12903z264), .I5 (nx12903z287)) ;
         defparam ix12903z17413.INIT = 64'h69F8921FCE213DC2;
    LUT6 ix42825z47621 (.O (px2828), .I0 (nx12903z459), .I1 (px2835), .I2 (
         nx12903z456), .I3 (nx12903z464), .I4 (nx12903z463), .I5 (nx12903z455)
         ) ;
         defparam ix42825z47621.INIT = 64'h648B6B741B5CB48B;
    LUT6 ix12903z40213 (.O (nx12903z455), .I0 (\p_key_samp(62)  ), .I1 (
         nx12903z258), .I2 (nx9305z10), .I3 (px3216), .I4 (px3010), .I5 (px2855)
         ) ;
         defparam ix12903z40213.INIT = 64'h9669699669969669;
    LUT6 ix12903z28745 (.O (nx12903z463), .I0 (\p_key_samp(30)  ), .I1 (
         nx12903z218), .I2 (px3483), .I3 (px3206), .I4 (px3006), .I5 (px2857)) ;
         defparam ix12903z28745.INIT = 64'h6996966996696996;
    LUT6 ix12903z28746 (.O (nx12903z464), .I0 (\p_key_samp(7)  ), .I1 (px3437), 
         .I2 (px3436), .I3 (px3197), .I4 (px3054), .I5 (px2832)) ;
         defparam ix12903z28746.INIT = 64'h6996966996696996;
    LUT6 ix12903z59873 (.O (px2832), .I0 (nx12903z394), .I1 (px2913), .I2 (
         px2912), .I3 (nx12903z409), .I4 (px2908), .I5 (px2906)) ;
         defparam ix12903z59873.INIT = 64'h996996592DD2E32C;
    LUT6 ix12903z28739 (.O (nx12903z456), .I0 (\p_key_samp(4)  ), .I1 (
         nx12903z457), .I2 (nx9305z5), .I3 (nx12903z111), .I4 (nx12903z352), .I5 (
         nx12903z458)) ;
         defparam ix12903z28739.INIT = 64'h6996966996696996;
    LUT6 ix12903z42384 (.O (nx12903z458), .I0 (px2879), .I1 (px2878), .I2 (
         px2877), .I3 (nx12903z440), .I4 (nx12903z445), .I5 (px2872)) ;
         defparam ix12903z42384.INIT = 64'hA97E439479069EE1;
    LUT6 ix43824z22735 (.O (px2836), .I0 (nx12903z264), .I1 (nx12903z287), .I2 (
         px2944), .I3 (px2942), .I4 (px2940), .I5 (px2928)) ;
         defparam ix43824z22735.INIT = 64'hDE35254AA4DC53A3;
    LUT6 ix12903z28742 (.O (nx12903z459), .I0 (\p_key_samp(39)  ), .I1 (
         nx12903z460), .I2 (nx9305z3), .I3 (nx12903z107), .I4 (nx12903z356), .I5 (
         nx12903z461)) ;
         defparam ix12903z28742.INIT = 64'h6996966996696996;
    LUT6 ix12903z34832 (.O (nx12903z461), .I0 (px2890), .I1 (nx12903z428), .I2 (
         px2884), .I3 (nx12903z434), .I4 (px2886), .I5 (px2887)) ;
         defparam ix12903z34832.INIT = 64'hDA8766347C96815E;
    LUT6 ix12903z40020 (.O (nx12903z213), .I0 (\p_key_samp(44)  ), .I1 (
         nx12903z214), .I2 (nx12903z6), .I3 (nx12903z94), .I4 (nx12903z131), .I5 (
         nx12903z215)) ;
         defparam ix12903z40020.INIT = 64'h9669699669969669;
    LUT6 ix12903z9103 (.O (nx12903z215), .I0 (px2866), .I1 (nx12903z217), .I2 (
         nx12903z257), .I3 (nx12903z260), .I4 (nx12903z303), .I5 (px2841)) ;
         defparam ix12903z9103.INIT = 64'h1A1DE3E4DC631DA2;
    LUT6 ix12903z40094 (.O (nx12903z303), .I0 (\p_key_samp(63)  ), .I1 (
         nx12903z304), .I2 (nx3326z8), .I3 (nx12903z99), .I4 (nx12903z135), .I5 (
         nx12903z305)) ;
         defparam ix12903z40094.INIT = 64'h9669699669969669;
    LUT6 ix12903z16381 (.O (nx12903z305), .I0 (nx12903z306), .I1 (nx12903z309), 
         .I2 (px2847), .I3 (px2846), .I4 (px2845), .I5 (px2844)) ;
         defparam ix12903z16381.INIT = 64'hA5C345795A3C39C6;
    LUT6 ix12903z28625 (.O (nx12903z309), .I0 (\p_key_samp(23)  ), .I1 (
         nx12903z310), .I2 (nx13298z29), .I3 (nx12903z58), .I4 (nx12903z139), .I5 (
         nx12903z311)) ;
         defparam ix12903z28625.INIT = 64'h6996966996696996;
    LUT6 ix12903z45967 (.O (nx12903z311), .I0 (px3053), .I1 (px3040), .I2 (
         nx12903z269), .I3 (px3034), .I4 (px3021), .I5 (nx12903z282)) ;
         defparam ix12903z45967.INIT = 64'h6B79148BD14EAD52;
    LUT6 ix12903z28622 (.O (nx12903z306), .I0 (\p_key_samp(53)  ), .I1 (
         nx12903z307), .I2 (nx13298z25), .I3 (nx12903z55), .I4 (nx12903z137), .I5 (
         nx12903z308)) ;
         defparam ix12903z28622.INIT = 64'h6996966996696996;
    LUT6 ix12903z40093 (.O (nx12903z308), .I0 (px2981), .I1 (nx12903z189), .I2 (
         nx12903z192), .I3 (px2972), .I4 (px2969), .I5 (px2966)) ;
         defparam ix12903z40093.INIT = 64'hD23C2DE4A5C69663;
    LUT6 ix12903z28585 (.O (nx12903z260), .I0 (\p_key_samp(20)  ), .I1 (
         nx12903z261), .I2 (nx3326z5), .I3 (nx12903z101), .I4 (nx12903z171), .I5 (
         nx12903z262)) ;
         defparam ix12903z28585.INIT = 64'h6996966996696996;
    LUT6 ix12903z59433 (.O (nx12903z262), .I0 (px2928), .I1 (nx12903z264), .I2 (
         px2942), .I3 (px2940), .I4 (nx12903z287), .I5 (px2944)) ;
         defparam ix12903z59433.INIT = 64'h619D3E611E72E11E;
    LUT6 ix12903z40057 (.O (nx12903z257), .I0 (\p_key_samp(46)  ), .I1 (
         nx12903z258), .I2 (nx9305z10), .I3 (px3216), .I4 (px3010), .I5 (px2855)
         ) ;
         defparam ix12903z40057.INIT = 64'h9669699669969669;
    LUT6 ix12903z18915 (.O (px2855), .I0 (px3056), .I1 (px3016), .I2 (
         nx12903z129), .I3 (px2984), .I4 (nx12903z185), .I5 (px2952)) ;
         defparam ix12903z18915.INIT = 64'h865A9E6CAD6643D1;
    LUT6 ix12903z28548 (.O (nx12903z217), .I0 (\p_key_samp(23)  ), .I1 (
         nx12903z218), .I2 (px3483), .I3 (px3206), .I4 (px3006), .I5 (px2857)) ;
         defparam ix12903z28548.INIT = 64'h6996966996696996;
    LUT6 ix12903z6613 (.O (px2857), .I0 (px2865), .I1 (nx12903z222), .I2 (
         nx12903z251), .I3 (px2860), .I4 (px2859), .I5 (px2858)) ;
         defparam ix12903z6613.INIT = 64'h53A5AF498C3B13E4;
    LUT5 ix12903z28579 (.O (nx12903z251), .I0 (\p_key_samp(15)  ), .I1 (
         nx12903z252), .I2 (nx32966z9), .I3 (nx12903z196), .I4 (nx12903z253)) ;
         defparam ix12903z28579.INIT = 32'h96696996;
    LUT6 ix12903z40315 (.O (nx12903z253), .I0 (px3015), .I1 (nx12903z133), .I2 (
         nx12903z164), .I3 (px3008), .I4 (px3005), .I5 (nx12903z169)) ;
         defparam ix12903z40315.INIT = 64'h64B309B6784B976C;
    LUT6 ix12903z28552 (.O (nx12903z222), .I0 (\p_key_samp(54)  ), .I1 (
         nx12903z223), .I2 (nx13298z50), .I3 (nx32966z7), .I4 (nx12903z200), .I5 (
         nx12903z224)) ;
         defparam ix12903z28552.INIT = 64'h6996966996696996;
    LUT6 ix12903z3517 (.O (nx12903z224), .I0 (px2939), .I1 (nx12903z226), .I2 (
         px2935), .I3 (px2934), .I4 (px2933), .I5 (nx12903z240)) ;
         defparam ix12903z3517.INIT = 64'h93A46E69589F07C9;
    LUT6 ix42825z36647 (.O (px2868), .I0 (nx61487z2), .I1 (px2926), .I2 (
         nx61487z5), .I3 (px2892), .I4 (nx61487z8), .I5 (px2870)) ;
         defparam ix42825z36647.INIT = 64'h66D178AE796989B0;
    LUT6 ix61487z51382 (.O (px2869), .I0 (nx61487z2), .I1 (px2926), .I2 (
         nx61487z5), .I3 (px2892), .I4 (nx61487z8), .I5 (px2870)) ;
         defparam ix61487z51382.INIT = 64'h51A8BA47ACF3C394;
    LUT6 ix42825z24686 (.O (px2871), .I0 (px2879), .I1 (px2878), .I2 (px2877), .I3 (
         nx12903z440), .I4 (nx12903z445), .I5 (px2872)) ;
         defparam ix42825z24686.INIT = 64'h3DC3605EC66C5AA5;
    LUT6 ix12903z28729 (.O (nx12903z445), .I0 (\p_key_samp(42)  ), .I1 (
         nx12903z446), .I2 (nx24265z26), .I3 (nx12903z22), .I4 (nx12903z232), .I5 (
         nx12903z447)) ;
         defparam ix12903z28729.INIT = 64'h6996966996696996;
    LUT6 ix12903z17291 (.O (nx12903z447), .I0 (px2924), .I1 (px2925), .I2 (
         px2921), .I3 (nx12903z403), .I4 (nx12903z406), .I5 (nx12903z399)) ;
         defparam ix12903z17291.INIT = 64'hC6ADCB12C9323CE5;
    LUT6 ix12903z40584 (.O (nx12903z440), .I0 (\p_key_samp(57)  ), .I1 (
         nx12903z441), .I2 (nx24265z37), .I3 (nx12903z20), .I4 (nx12903z235), .I5 (
         nx12903z442)) ;
         defparam ix12903z40584.INIT = 64'h9669699669969669;
    LUT6 ix12903z35311 (.O (nx12903z442), .I0 (nx12903z342), .I1 (px3076), .I2 (
         nx12903z345), .I3 (px3059), .I4 (px3089), .I5 (nx12903z340)) ;
         defparam ix12903z35311.INIT = 64'hA6AD78D16E92834D;
    LUT6 ix61487z39824 (.O (nx61487z8), .I0 (\p_key_samp(14)  ), .I1 (px3521), .I2 (
         px3506), .I3 (px3313), .I4 (px3090), .I5 (px2881)) ;
         defparam ix61487z39824.INIT = 64'h9669699669969669;
    LUT6 ix61487z28180 (.O (px2881), .I0 (px2890), .I1 (nx12903z428), .I2 (
         px2887), .I3 (px2886), .I4 (px2884), .I5 (nx12903z434)) ;
         defparam ix61487z28180.INIT = 64'h7289C519975C68EB;
    LUT6 ix12903z28719 (.O (nx12903z434), .I0 (\p_key_samp(13)  ), .I1 (
         nx12903z435), .I2 (nx7312z12), .I3 (nx12903z36), .I4 (nx12903z363), .I5 (
         nx12903z436)) ;
         defparam ix12903z28719.INIT = 64'h6996966996696996;
    LUT6 ix12903z59393 (.O (nx12903z436), .I0 (nx12903z226), .I1 (px2934), .I2 (
         px2935), .I3 (px2933), .I4 (nx12903z240), .I5 (px2939)) ;
         defparam ix12903z59393.INIT = 64'hE1961EB19C4BE166;
    LUT6 ix42825z52111 (.O (px2885), .I0 (px2925), .I1 (px2924), .I2 (
         nx12903z399), .I3 (px2921), .I4 (nx12903z403), .I5 (nx12903z406)) ;
         defparam ix42825z52111.INIT = 64'h6336E89C966CC659;
    LUT6 ix12903z40190 (.O (nx12903z428), .I0 (\p_key_samp(22)  ), .I1 (
         nx12903z429), .I2 (nx7312z17), .I3 (nx12903z31), .I4 (nx12903z360), .I5 (
         nx12903z430)) ;
         defparam ix12903z40190.INIT = 64'h9669699669969669;
    LUT6 ix12903z26957 (.O (nx12903z430), .I0 (px2999), .I1 (nx12903z295), .I2 (
         px2996), .I3 (nx12903z292), .I4 (nx12903z298), .I5 (px2986)) ;
         defparam ix12903z26957.INIT = 64'hD0C3BC0F2D5A62B5;
    LUT6 ix42825z47510 (.O (px2891), .I0 (px3015), .I1 (nx12903z133), .I2 (
         nx12903z164), .I3 (px3008), .I4 (px3005), .I5 (nx12903z169)) ;
         defparam ix42825z47510.INIT = 64'h3D924B69C29DB463;
    LUT6 ix42825z29335 (.O (px2893), .I0 (nx12903z334), .I1 (nx12903z346), .I2 (
         px2898), .I3 (px2897), .I4 (px2896), .I5 (px2894)) ;
         defparam ix42825z29335.INIT = 64'hC653996D953A6CC2;
    LUT6 ix42825z27162 (.O (px2895), .I0 (px2925), .I1 (px2924), .I2 (
         nx12903z399), .I3 (px2921), .I4 (nx12903z403), .I5 (nx12903z406)) ;
         defparam ix42825z27162.INIT = 64'hC36C9659B97A6494;
    LUT6 ix42825z28921 (.O (px2899), .I0 (px3053), .I1 (px3040), .I2 (
         nx12903z269), .I3 (px3034), .I4 (px3021), .I5 (nx12903z282)) ;
         defparam ix42825z28921.INIT = 64'h521A8DE2B8D76B94;
    LUT6 ix12903z28651 (.O (nx12903z346), .I0 (\p_key_samp(34)  ), .I1 (
         nx12903z347), .I2 (nx13298z65), .I3 (nx12903z77), .I4 (nx12903z279), .I5 (
         nx12903z348)) ;
         defparam ix12903z28651.INIT = 64'h6996966996696996;
    LUT6 ix12903z55293 (.O (nx12903z348), .I0 (px2963), .I1 (nx12903z350), .I2 (
         px2959), .I3 (nx12903z354), .I4 (nx12903z365), .I5 (nx12903z366)) ;
         defparam ix12903z55293.INIT = 64'h46ABA1D9619ED1A6;
    LUT6 ix12903z28642 (.O (nx12903z334), .I0 (\p_key_samp(52)  ), .I1 (
         nx12903z335), .I2 (nx13298z62), .I3 (nx12903z79), .I4 (nx12903z277), .I5 (
         nx12903z336)) ;
         defparam ix12903z28642.INIT = 64'h6996966996696996;
    LUT6 ix12903z59860 (.O (nx12903z336), .I0 (px3089), .I1 (px3076), .I2 (
         px3059), .I3 (nx12903z340), .I4 (nx12903z342), .I5 (nx12903z345)) ;
         defparam ix12903z59860.INIT = 64'hE79A54291675E386;
    LUT6 ix61487z39822 (.O (nx61487z5), .I0 (\p_key_samp(31)  ), .I1 (nx61487z6)
         , .I2 (nx11304z6), .I3 (nx12903z88), .I4 (nx12903z344), .I5 (
         nx12903z393)) ;
         defparam ix61487z39822.INIT = 64'h9669699669969669;
    LUT6 ix12903z48834 (.O (nx12903z393), .I0 (nx12903z394), .I1 (px2913), .I2 (
         px2912), .I3 (nx12903z409), .I4 (px2908), .I5 (px2906)) ;
         defparam ix12903z48834.INIT = 64'hE93E1EB86641B847;
    LUT6 ix12903z38230 (.O (px2907), .I0 (px2999), .I1 (px2996), .I2 (
         nx12903z292), .I3 (nx12903z295), .I4 (nx12903z298), .I5 (px2986)) ;
         defparam ix12903z38230.INIT = 64'h2D90D36E533E8E94;
    LUT6 ix56500z27230 (.O (px2909), .I0 (px2969), .I1 (px2972), .I2 (px2981), .I3 (
         nx12903z189), .I4 (nx12903z192), .I5 (px2966)) ;
         defparam ix56500z27230.INIT = 64'h6D305AC75AC6653C;
    LUT6 ix12903z40177 (.O (nx12903z409), .I0 (\p_key_samp(47)  ), .I1 (
         nx12903z410), .I2 (nx13298z46), .I3 (nx12903z46), .I4 (nx12903z246), .I5 (
         nx12903z411)) ;
         defparam ix12903z40177.INIT = 64'h9669699669969669;
    LUT6 ix12903z44116 (.O (nx12903z411), .I0 (px2963), .I1 (nx12903z350), .I2 (
         px2959), .I3 (nx12903z354), .I4 (nx12903z365), .I5 (nx12903z366)) ;
         defparam ix12903z44116.INIT = 64'h87D2C996782DA5CA;
    LUT6 ix12903z57629 (.O (px2914), .I0 (px2939), .I1 (nx12903z226), .I2 (
         px2935), .I3 (px2934), .I4 (px2933), .I5 (nx12903z240)) ;
         defparam ix12903z57629.INIT = 64'h6B8324F839D4DA65;
    LUT6 ix12903z28690 (.O (nx12903z394), .I0 (\p_key_samp(4)  ), .I1 (
         nx12903z395), .I2 (nx13298z39), .I3 (nx12903z41), .I4 (nx12903z244), .I5 (
         nx12903z396)) ;
         defparam ix12903z28690.INIT = 64'h6996966996696996;
    LUT6 ix12903z28744 (.O (nx12903z396), .I0 (px2925), .I1 (px2924), .I2 (
         nx12903z399), .I3 (px2921), .I4 (nx12903z403), .I5 (nx12903z406)) ;
         defparam ix12903z28744.INIT = 64'h39C68E35873969CA;
    LUT6 ix12903z40176 (.O (nx12903z406), .I0 (\p_key_samp(33)  ), .I1 (px3714)
         , .I2 (px3705), .I3 (px3460), .I4 (px3232), .I5 (px2973)) ;
         defparam ix12903z40176.INIT = 64'h9669699669969669;
    LUT6 ix12903z28698 (.O (nx12903z403), .I0 (\p_key_samp(3)  ), .I1 (
         nx12903z404), .I2 (nx24265z33), .I3 (nx337z4), .I4 (nx12903z145), .I5 (
         nx12903z405)) ;
         defparam ix12903z28698.INIT = 64'h6996966996696996;
    LUT6 ix12903z32015 (.O (nx12903z405), .I0 (nx12903z272), .I1 (nx12903z273), 
         .I2 (nx12903z274), .I3 (nx12903z275), .I4 (nx12903z276), .I5 (
         nx12903z278)) ;
         defparam ix12903z32015.INIT = 64'hAC5613E6C93A7689;
    (* HLUTNM = "LUT62_1_29" *)
    LUT5 ix45810z28362 (.O (nx45810z19), .I0 (\plaintext(16)  ), .I1 (nx34235z28
         ), .I2 (nx24265z33), .I3 (nx337z4), .I4 (nx12903z145)) ;
         defparam ix45810z28362.INIT = 32'h96696996;
    LUT6 ix12903z28693 (.O (nx12903z399), .I0 (\p_key_samp(60)  ), .I1 (
         nx12903z400), .I2 (nx24265z31), .I3 (nx337z6), .I4 (nx12903z147), .I5 (
         nx12903z401)) ;
         defparam ix12903z28693.INIT = 64'h6996966996696996;
    LUT6 ix12903z28889 (.O (nx12903z401), .I0 (nx12903z357), .I1 (nx12903z359), 
         .I2 (nx12903z362), .I3 (nx12903z361), .I4 (nx12903z358), .I5 (
         nx12903z364)) ;
         defparam ix12903z28889.INIT = 64'h7AE18D93934C68F4;
    LUT6 ix42825z16438 (.O (px2927), .I0 (nx12903z264), .I1 (nx12903z287), .I2 (
         px2944), .I3 (px2942), .I4 (px2940), .I5 (px2928)) ;
         defparam ix42825z16438.INIT = 64'h39ACC66BA5323A95;
    LUT6 ix42825z20988 (.O (px2929), .I0 (px2939), .I1 (nx12903z226), .I2 (
         px2935), .I3 (px2934), .I4 (px2933), .I5 (nx12903z240)) ;
         defparam ix42825z20988.INIT = 64'h16EABC4B334D4CB4;
    LUT6 ix12903z28568 (.O (nx12903z240), .I0 (\p_key_samp(27)  ), .I1 (
         nx12903z241), .I2 (nx24265z23), .I3 (nx4319z3), .I4 (nx12903z160), .I5 (
         nx12903z242)) ;
         defparam ix12903z28568.INIT = 64'h6996966996696996;
    LUT6 ix12903z16541 (.O (nx12903z242), .I0 (nx12903z243), .I1 (nx12903z245), 
         .I2 (nx12903z247), .I3 (nx12903z248), .I4 (nx12903z249), .I5 (
         nx12903z250)) ;
         defparam ix12903z16541.INIT = 64'hC63AC5A5C35A3A99;
    (* HLUTNM = "LUT62_1_22" *)
    LUT5 ix44815z39841 (.O (nx44815z23), .I0 (\plaintext(10)  ), .I1 (nx29253z10
         ), .I2 (nx24265z23), .I3 (nx4319z3), .I4 (nx12903z160)) ;
         defparam ix44815z39841.INIT = 32'h69969669;
    LUT6 ix12903z40030 (.O (nx12903z226), .I0 (\p_key_samp(44)  ), .I1 (
         nx12903z227), .I2 (nx24265z20), .I3 (nx4319z5), .I4 (nx12903z163), .I5 (
         nx12903z228)) ;
         defparam ix12903z40030.INIT = 64'h9669699669969669;
    LUT6 ix12903z44900 (.O (nx12903z228), .I0 (nx12903z229), .I1 (nx12903z230), 
         .I2 (nx12903z231), .I3 (nx12903z233), .I4 (nx12903z234), .I5 (
         nx12903z236)) ;
         defparam ix12903z44900.INIT = 64'h9A59536C65B1A96C;
    (* HLUTNM = "LUT62_1_21" *)
    LUT5 ix44815z39838 (.O (nx44815z20), .I0 (\plaintext(18)  ), .I1 (nx29253z8)
         , .I2 (nx24265z20), .I3 (nx4319z5), .I4 (nx12903z163)) ;
         defparam ix44815z39838.INIT = 32'h69969669;
    LUT6 ix42825z45769 (.O (px2941), .I0 (px3005), .I1 (nx12903z133), .I2 (
         nx12903z169), .I3 (px3008), .I4 (nx12903z164), .I5 (px3015)) ;
         defparam ix42825z45769.INIT = 64'hB178468F4E87AD70;
    LUT6 ix42825z54975 (.O (px2943), .I0 (px2969), .I1 (nx12903z192), .I2 (
         nx12903z189), .I3 (px2981), .I4 (px2972), .I5 (px2966)) ;
         defparam ix42825z54975.INIT = 64'hD829A5D62DD2D16A;
    LUT6 ix42825z39804 (.O (px2945), .I0 (px2959), .I1 (nx12903z366), .I2 (
         nx12903z350), .I3 (px2963), .I4 (nx12903z365), .I5 (nx12903z354)) ;
         defparam ix42825z39804.INIT = 64'hC57A3CC36A92962D;
    LUT6 ix12903z28606 (.O (nx12903z287), .I0 (\p_key_samp(19)  ), .I1 (
         nx12903z288), .I2 (nx13298z9), .I3 (nx35956z6), .I4 (nx12903z177), .I5 (
         nx12903z289)) ;
         defparam ix12903z28606.INIT = 64'h6996966996696996;
    LUT6 ix12903z39408 (.O (nx12903z289), .I0 (px2999), .I1 (px2996), .I2 (
         nx12903z292), .I3 (nx12903z295), .I4 (nx12903z298), .I5 (px2986)) ;
         defparam ix12903z39408.INIT = 64'h56969AA56D9293C6;
    LUT6 ix12903z28589 (.O (nx12903z264), .I0 (\p_key_samp(9)  ), .I1 (
         nx12903z265), .I2 (nx13298z5), .I3 (nx35956z4), .I4 (nx12903z175), .I5 (
         nx12903z266)) ;
         defparam ix12903z28589.INIT = 64'h6996966996696996;
    LUT6 ix12903z43678 (.O (nx12903z266), .I0 (px3053), .I1 (px3040), .I2 (
         nx12903z269), .I3 (px3034), .I4 (px3021), .I5 (nx12903z282)) ;
         defparam ix12903z43678.INIT = 64'h16E9D72E8B72A485;
    LUT6 ix61487z28345 (.O (nx61487z2), .I0 (\p_key_samp(5)  ), .I1 (nx61487z3)
         , .I2 (nx11304z3), .I3 (nx12903z4), .I4 (nx12903z13), .I5 (nx12903z126)
         ) ;
         defparam ix61487z28345.INIT = 64'h6996966996696996;
    LUT6 ix12903z32744 (.O (nx12903z126), .I0 (px3056), .I1 (px3016), .I2 (
         nx12903z129), .I3 (px2984), .I4 (nx12903z185), .I5 (px2952)) ;
         defparam ix12903z32744.INIT = 64'h9B5CC48B64D37A49;
    LUT6 ix42825z19746 (.O (px2953), .I0 (px2963), .I1 (nx12903z350), .I2 (
         px2959), .I3 (nx12903z354), .I4 (nx12903z365), .I5 (nx12903z366)) ;
         defparam ix42825z19746.INIT = 64'h2BE1B41E3C5647A9;
    LUT6 ix12903z28670 (.O (nx12903z366), .I0 (\p_key_samp(4)  ), .I1 (px3636), 
         .I2 (px3635), .I3 (px3436), .I4 (px3197), .I5 (px3054)) ;
         defparam ix12903z28670.INIT = 64'h6996966996696996;
    LUT6 ix12903z28669 (.O (nx12903z365), .I0 (\p_key_samp(30)  ), .I1 (
         nx12903z165), .I2 (nx36230z11), .I3 (nx9305z10), .I4 (px3216), .I5 (
         px3010)) ;
         defparam ix12903z28669.INIT = 64'h6996966996696996;
    LUT6 ix12903z40133 (.O (nx12903z354), .I0 (\p_key_samp(7)  ), .I1 (
         nx12903z355), .I2 (nx36230z3), .I3 (nx9305z3), .I4 (nx12903z107), .I5 (
         nx12903z356)) ;
         defparam ix12903z40133.INIT = 64'h9669699669969669;
    LUT6 ix12903z28058 (.O (nx12903z356), .I0 (nx12903z357), .I1 (nx12903z358), 
         .I2 (nx12903z359), .I3 (nx12903z361), .I4 (nx12903z362), .I5 (
         nx12903z364)) ;
         defparam ix12903z28058.INIT = 64'h7AC4C193AD92673C;
    (* HLUTNM = "LUT62_1_14" *)
    LUT5 ix43820z28351 (.O (nx43820z9), .I0 (\plaintext(12)  ), .I1 (nx37232z4)
         , .I2 (nx36230z3), .I3 (nx9305z3), .I4 (nx12903z107)) ;
         defparam ix43820z28351.INIT = 32'h96696996;
    LUT6 ix12903z28654 (.O (nx12903z350), .I0 (\p_key_samp(37)  ), .I1 (
         nx12903z351), .I2 (nx36230z5), .I3 (nx9305z5), .I4 (nx12903z111), .I5 (
         nx12903z352)) ;
         defparam ix12903z28654.INIT = 64'h6996966996696996;
    LUT6 ix12903z35284 (.O (nx12903z352), .I0 (nx12903z231), .I1 (nx12903z236), 
         .I2 (nx12903z233), .I3 (nx12903z229), .I4 (nx12903z230), .I5 (
         nx12903z234)) ;
         defparam ix12903z35284.INIT = 64'hA5D97C86591A8379;
    (* HLUTNM = "LUT62_1_15" *)
    LUT5 ix43820z28355 (.O (nx43820z14), .I0 (\plaintext(20)  ), .I1 (nx37232z6)
         , .I2 (nx36230z5), .I3 (nx9305z5), .I4 (nx12903z111)) ;
         defparam ix43820z28355.INIT = 32'h96696996;
    LUT6 ix12903z39998 (.O (nx12903z185), .I0 (\p_key_samp(60)  ), .I1 (
         nx12903z186), .I2 (nx13298z72), .I3 (nx12903z8), .I4 (nx12903z61), .I5 (
         nx12903z187)) ;
         defparam ix12903z39998.INIT = 64'h9669699669969669;
    LUT6 ix12903z62982 (.O (nx12903z187), .I0 (px2981), .I1 (nx12903z189), .I2 (
         nx12903z192), .I3 (px2972), .I4 (px2969), .I5 (px2966)) ;
         defparam ix12903z62982.INIT = 64'h99A56E52139CF02F;
    LUT6 ix44815z20187 (.O (px2967), .I0 (nx12903z357), .I1 (nx12903z358), .I2 (
         nx12903z359), .I3 (nx12903z361), .I4 (nx12903z364), .I5 (nx12903z362)
         ) ;
         defparam ix44815z20187.INIT = 64'hC9833CE6235E49B5;
    (* HLUTNM = "LUT62_1_19" *)
    LUT5 ix44815z28347 (.O (nx44815z4), .I0 (\plaintext(26)  ), .I1 (nx45210z2)
         , .I2 (px3716), .I3 (px3454), .I4 (px3226)) ;
         defparam ix44815z28347.INIT = 32'h96696996;
    LUT6 ix12903z12983 (.O (px2970), .I0 (nx12903z272), .I1 (nx12903z273), .I2 (
         nx12903z274), .I3 (nx12903z275), .I4 (nx12903z276), .I5 (nx12903z278)
         ) ;
         defparam ix12903z12983.INIT = 64'h964AB6935AB42C6D;
    (* HLUTNM = "LUT62_1_20" *)
    LUT5 ix44815z39828 (.O (nx44815z10), .I0 (\plaintext(34)  ), .I1 (nx41222z2)
         , .I2 (px3688), .I3 (px3448), .I4 (px3229)) ;
         defparam ix44815z39828.INIT = 32'h69969669;
    LUT6 ix12903z33035 (.O (px2973), .I0 (nx12903z152), .I1 (nx12903z150), .I2 (
         nx12903z136), .I3 (nx12903z140), .I4 (nx12903z138), .I5 (nx12903z154)
         ) ;
         defparam ix12903z33035.INIT = 64'h2D96C33C926A7AC5;
    (* HLUTNM = "LUT62_1_26" *)
    LUT5 ix44819z39829 (.O (nx44819z11), .I0 (\plaintext(58)  ), .I1 (nx34235z18
         ), .I2 (px3705), .I3 (px3460), .I4 (px3232)) ;
         defparam ix44819z39829.INIT = 32'h69969669;
    LUT6 ix12903z28529 (.O (nx12903z192), .I0 (\p_key_samp(41)  ), .I1 (
         nx12903z193), .I2 (nx7313z10), .I3 (nx7312z7), .I4 (nx12903z63), .I5 (
         nx12903z194)) ;
         defparam ix12903z28529.INIT = 64'h6996966996696996;
    LUT6 ix12903z37056 (.O (nx12903z194), .I0 (nx12903z195), .I1 (nx12903z197), 
         .I2 (nx12903z199), .I3 (nx12903z201), .I4 (nx12903z203), .I5 (
         nx12903z205)) ;
         defparam ix12903z37056.INIT = 64'h55E9691DC3168AE3;
    (* HLUTNM = "LUT62_1_25" *)
    LUT5 ix44819z39826 (.O (nx44819z8), .I0 (\plaintext(50)  ), .I1 (nx34235z13)
         , .I2 (nx7313z10), .I3 (nx7312z7), .I4 (nx12903z63)) ;
         defparam ix44819z39826.INIT = 32'h69969669;
    LUT6 ix12903z40001 (.O (nx12903z189), .I0 (\p_key_samp(26)  ), .I1 (
         nx12903z190), .I2 (nx7313z4), .I3 (nx7312z3), .I4 (nx12903z65), .I5 (
         nx12903z191)) ;
         defparam ix12903z40001.INIT = 64'h9669699669969669;
    LUT6 ix12903z7363 (.O (nx12903z191), .I0 (nx12903z182), .I1 (nx12903z176), .I2 (
         nx12903z180), .I3 (nx12903z174), .I4 (nx12903z178), .I5 (nx12903z172)
         ) ;
         defparam ix12903z7363.INIT = 64'h31C37827ED1C16E9;
    (* HLUTNM = "LUT62_1_23" *)
    LUT5 ix44819z28348 (.O (nx44819z5), .I0 (\plaintext(42)  ), .I1 (nx34235z15)
         , .I2 (nx7313z4), .I3 (nx7312z3), .I4 (nx12903z65)) ;
         defparam ix44819z28348.INIT = 32'h96696996;
    LUT6 ix44819z43166 (.O (px2982), .I0 (nx12903z104), .I1 (nx12903z60), .I2 (
         nx12903z14), .I3 (nx12903z115), .I4 (nx12903z93), .I5 (nx12903z82)) ;
         defparam ix44819z43166.INIT = 64'hA9D45C0B7666A36C;
    (* HLUTNM = "LUT62_1_24" *)
    LUT5 ix44819z28359 (.O (nx44819z16), .I0 (plaintext[6]), .I1 (nx44209z2), .I2 (
         px3702), .I3 (px3451), .I4 (px3235)) ;
         defparam ix44819z28359.INIT = 32'h96696996;
    LUT6 ix12903z40616 (.O (px2985), .I0 (px2999), .I1 (px2996), .I2 (
         nx12903z292), .I3 (nx12903z295), .I4 (nx12903z298), .I5 (px2986)) ;
         defparam ix12903z40616.INIT = 64'h4B3536E8D4CA9837;
    LUT6 ix45810z7061 (.O (px2987), .I0 (nx12903z243), .I1 (nx12903z248), .I2 (
         nx12903z249), .I3 (nx12903z245), .I4 (nx12903z250), .I5 (nx12903z247)
         ) ;
         defparam ix45810z7061.INIT = 64'h1497E36CE9991666;
    (* HLUTNM = "LUT62_1_28" *)
    LUT5 ix45810z28356 (.O (nx45810z13), .I0 (\plaintext(24)  ), .I1 (nx39226z17
         ), .I2 (px3657), .I3 (px3410), .I4 (px3261)) ;
         defparam ix45810z28356.INIT = 32'h96696996;
    LUT6 ix12903z40091 (.O (nx12903z298), .I0 (\p_key_samp(18)  ), .I1 (
         nx12903z299), .I2 (nx24265z12), .I3 (nx5318z9), .I4 (nx12903z51), .I5 (
         nx12903z300)) ;
         defparam ix12903z40091.INIT = 64'h9669699669969669;
    LUT6 ix12903z29648 (.O (nx12903z300), .I0 (nx12903z136), .I1 (nx12903z138), 
         .I2 (nx12903z140), .I3 (nx12903z150), .I4 (nx12903z152), .I5 (
         nx12903z154)) ;
         defparam ix12903z29648.INIT = 64'hCB3E58942C696D9C;
    (* HLUTNM = "LUT62_1_31" *)
    LUT5 ix45814z39829 (.O (nx45814z11), .I0 (\plaintext(40)  ), .I1 (nx39226z7)
         , .I2 (nx24265z12), .I3 (nx5318z9), .I4 (nx12903z51)) ;
         defparam ix45814z39829.INIT = 32'h69969669;
    LUT6 ix12903z28613 (.O (nx12903z295), .I0 (\p_key_samp(11)  ), .I1 (
         nx12903z296), .I2 (nx27254z2), .I3 (px3536), .I4 (px3330), .I5 (px3136)
         ) ;
         defparam ix12903z28613.INIT = 64'h6996966996696996;
    LUT6 ix12903z28609 (.O (nx12903z292), .I0 (\p_key_samp(36)  ), .I1 (
         nx12903z293), .I2 (nx24265z7), .I3 (nx5318z6), .I4 (nx12903z27), .I5 (
         nx12903z294)) ;
         defparam ix12903z28609.INIT = 64'h6996966996696996;
    LUT6 ix12903z29449 (.O (nx12903z294), .I0 (nx12903z201), .I1 (nx12903z205), 
         .I2 (nx12903z203), .I3 (nx12903z199), .I4 (nx12903z195), .I5 (
         nx12903z197)) ;
         defparam ix12903z29449.INIT = 64'h49DAB32986316CDB;
    (* HLUTNM = "LUT62_1_30" *)
    LUT5 ix45814z28351 (.O (nx45814z8), .I0 (\plaintext(48)  ), .I1 (nx39226z4)
         , .I2 (nx24265z7), .I3 (nx5318z6), .I4 (nx12903z27)) ;
         defparam ix45814z28351.INIT = 32'h96696996;
    LUT6 ix12903z39680 (.O (px2997), .I0 (nx12903z234), .I1 (nx12903z231), .I2 (
         nx12903z229), .I3 (nx12903z233), .I4 (nx12903z236), .I5 (nx12903z230)
         ) ;
         defparam ix12903z39680.INIT = 64'h3C276BD2A39C9463;
    (* HLUTNM = "LUT62_1_27" *)
    LUT5 ix45810z28349 (.O (nx45810z6), .I0 (\plaintext(32)  ), .I1 (nx39226z15)
         , .I2 (px3665), .I3 (px3421), .I4 (px3278)) ;
         defparam ix45810z28349.INIT = 32'h96696996;
    LUT6 ix12903z39945 (.O (nx12903z129), .I0 (\p_key_samp(43)  ), .I1 (
         nx12903z130), .I2 (nx13298z76), .I3 (nx12903z6), .I4 (nx12903z94), .I5 (
         nx12903z131)) ;
         defparam ix12903z39945.INIT = 64'h9669699669969669;
    LUT6 ix12903z56364 (.O (nx12903z131), .I0 (px3015), .I1 (nx12903z133), .I2 (
         nx12903z164), .I3 (px3008), .I4 (px3005), .I5 (nx12903z169)) ;
         defparam ix12903z56364.INIT = 64'hBC0626751CF3D68A;
    LUT6 ix12903z28508 (.O (nx12903z169), .I0 (\p_key_samp(53)  ), .I1 (
         nx12903z170), .I2 (nx13298z15), .I3 (nx3326z5), .I4 (nx12903z101), .I5 (
         nx12903z171)) ;
         defparam ix12903z28508.INIT = 64'h6996966996696996;
    (* HLUTNM = "LUT62_1_10" *)
    LUT5 ix43816z28348 (.O (nx43816z5), .I0 (\plaintext(54)  ), .I1 (nx34235z34)
         , .I2 (nx13298z15), .I3 (nx3326z5), .I4 (nx12903z101)) ;
         defparam ix43816z28348.INIT = 32'h96696996;
    LUT6 ix12903z55285 (.O (nx12903z171), .I0 (nx12903z172), .I1 (nx12903z174), 
         .I2 (nx12903z176), .I3 (nx12903z178), .I4 (nx12903z180), .I5 (
         nx12903z182)) ;
         defparam ix12903z55285.INIT = 64'h962E2BD139D2D22D;
    LUT6 ix12903z64386 (.O (px3006), .I0 (nx12903z197), .I1 (nx12903z199), .I2 (
         nx12903z195), .I3 (nx12903z205), .I4 (nx12903z203), .I5 (nx12903z201)
         ) ;
         defparam ix12903z64386.INIT = 64'h31DCC827CAA5F592;
    (* HLUTNM = "LUT62_1_1" *)
    LUT5 ix32966z39819 (.O (px3007), .I0 (plaintext[2]), .I1 (nx40221z2), .I2 (
         px3674), .I3 (px3483), .I4 (px3206)) ;
         defparam ix32966z39819.INIT = 32'h69969669;
    LUT6 ix12903z28505 (.O (nx12903z164), .I0 (\p_key_samp(14)  ), .I1 (
         nx12903z165), .I2 (nx36230z11), .I3 (nx9305z10), .I4 (px3216), .I5 (
         px3010)) ;
         defparam ix12903z28505.INIT = 64'h6996966996696996;
    LUT6 ix12903z24550 (.O (px3010), .I0 (nx12903z14), .I1 (nx12903z60), .I2 (
         nx12903z82), .I3 (nx12903z93), .I4 (nx12903z104), .I5 (nx12903z115)) ;
         defparam ix12903z24550.INIT = 64'h7C2997F816CE5A21;
    (* HLUTNM = "LUT62_1_12" *)
    LUT5 ix43816z39836 (.O (nx43816z22), .I0 (\plaintext(62)  ), .I1 (nx37232z13
         ), .I2 (nx36230z11), .I3 (nx9305z10), .I4 (px3216)) ;
         defparam ix43816z39836.INIT = 32'h69969669;
    LUT6 ix12903z39948 (.O (nx12903z133), .I0 (\p_key_samp(31)  ), .I1 (
         nx12903z134), .I2 (nx13298z13), .I3 (nx3326z8), .I4 (nx12903z99), .I5 (
         nx12903z135)) ;
         defparam ix12903z39948.INIT = 64'h9669699669969669;
    LUT6 ix12903z15215 (.O (nx12903z135), .I0 (nx12903z136), .I1 (nx12903z138), 
         .I2 (nx12903z140), .I3 (nx12903z150), .I4 (nx12903z152), .I5 (
         nx12903z154)) ;
         defparam ix12903z15215.INIT = 64'h6A8B963CCA3535CA;
    (* HLUTNM = "LUT62_1_11" *)
    LUT5 ix43816z39827 (.O (nx43816z9), .I0 (\plaintext(46)  ), .I1 (nx34235z37)
         , .I2 (nx13298z13), .I3 (nx3326z8), .I4 (nx12903z99)) ;
         defparam ix43816z39827.INIT = 32'h69969669;
    LUT6 ix33963z29451 (.O (px3017), .I0 (px3053), .I1 (px3040), .I2 (
         nx12903z269), .I3 (px3034), .I4 (px3021), .I5 (nx12903z282)) ;
         defparam ix33963z29451.INIT = 64'h857AB147E2146DE9;
    LUT6 ix12903z28603 (.O (nx12903z282), .I0 (\p_key_samp(62)  ), .I1 (
         nx12903z283), .I2 (nx15291z38), .I3 (nx13298z70), .I4 (nx12903z123), .I5 (
         nx12903z284)) ;
         defparam ix12903z28603.INIT = 64'h6996966996696996;
    LUT6 ix12903z51284 (.O (nx12903z284), .I0 (nx12903z60), .I1 (nx12903z104), .I2 (
         nx12903z93), .I3 (nx12903z14), .I4 (nx12903z82), .I5 (nx12903z115)) ;
         defparam ix12903z51284.INIT = 64'hB6581DE66993C22D;
    (* HLUTNM = "LUT62_1_16" *)
    LUT5 ix43824z28350 (.O (nx43824z8), .I0 (\plaintext(44)  ), .I1 (nx36228z4)
         , .I2 (nx15291z38), .I3 (nx13298z70), .I4 (nx12903z123)) ;
         defparam ix43824z28350.INIT = 32'h96696996;
    LUT6 ix42825z22757 (.O (px3022), .I0 (nx12903z136), .I1 (nx12903z138), .I2 (
         nx12903z140), .I3 (nx12903z150), .I4 (nx12903z152), .I5 (nx12903z154)
         ) ;
         defparam ix42825z22757.INIT = 64'h532CAC798DD153A6;
    LUT6 ix12903z39970 (.O (nx12903z154), .I0 (\p_plaintext(63)  ), .I1 (
         \p_key_samp(14)  ), .I2 (nx29253z2), .I3 (px3565), .I4 (px3359), .I5 (
         px3119)) ;
         defparam ix12903z39970.INIT = 64'h9669699669969669;
    LUT6 ix12903z28493 (.O (nx12903z152), .I0 (p_nbus_plaintext[63]), .I1 (
         \p_key_samp(47)  ), .I2 (nx63157z2), .I3 (px3724), .I4 (px3504), .I5 (
         px3281)) ;
         defparam ix12903z28493.INIT = 64'h6996966996696996;
    LUT6 ix12903z28491 (.O (nx12903z150), .I0 (\p_plaintext(37)  ), .I1 (
         \p_key_samp(53)  ), .I2 (px3745), .I3 (px3514), .I4 (px3315), .I5 (
         px3092)) ;
         defparam ix12903z28491.INIT = 64'h6996966996696996;
    LUT6 ix12903z28480 (.O (nx12903z140), .I0 (\plaintext(29)  ), .I1 (
         \p_key_samp(38)  ), .I2 (nx23267z2), .I3 (px3511), .I4 (px3321), .I5 (
         px3095)) ;
         defparam ix12903z28480.INIT = 64'h6996966996696996;
    LUT6 ix12903z28478 (.O (nx12903z138), .I0 (\plaintext(13)  ), .I1 (
         \p_key_samp(20)  ), .I2 (nx15291z29), .I3 (nx13298z29), .I4 (nx12903z58
         ), .I5 (nx12903z139)) ;
         defparam ix12903z28478.INIT = 64'h6996966996696996;
    LUT6 ix12903z7547 (.O (nx12903z139), .I0 (nx12903z117), .I1 (nx12903z118), .I2 (
         nx12903z119), .I3 (nx12903z120), .I4 (nx12903z122), .I5 (nx12903z124)
         ) ;
         defparam ix12903z7547.INIT = 64'h42E13C87B96E17D2;
    (* HLUTNM = "LUT62_1_51" *)
    LUT4 ix43816z28358 (.O (nx43816z17), .I0 (\plaintext(13)  ), .I1 (nx15291z29
         ), .I2 (nx13298z29), .I3 (nx12903z58)) ;
         defparam ix43816z28358.INIT = 16'h6996;
    LUT6 ix12903z28476 (.O (nx12903z136), .I0 (\plaintext(21)  ), .I1 (
         \p_key_samp(21)  ), .I2 (nx15291z32), .I3 (nx13298z25), .I4 (nx12903z55
         ), .I5 (nx12903z137)) ;
         defparam ix12903z28476.INIT = 64'h6996966996696996;
    LUT6 ix12903z28736 (.O (nx12903z137), .I0 (nx12903z62), .I1 (nx12903z64), .I2 (
         nx12903z66), .I3 (nx12903z68), .I4 (nx12903z70), .I5 (nx12903z80)) ;
         defparam ix12903z28736.INIT = 64'h69C6A56395A36A99;
    (* HLUTNM = "LUT62_1_50" *)
    LUT4 ix43816z28355 (.O (nx43816z12), .I0 (\plaintext(21)  ), .I1 (nx15291z32
         ), .I2 (nx13298z25), .I3 (nx12903z55)) ;
         defparam ix43816z28355.INIT = 16'h6996;
    (* HLUTNM = "LUT62_1_17" *)
    LUT5 ix43824z28358 (.O (nx43824z16), .I0 (\plaintext(60)  ), .I1 (nx36228z10
         ), .I2 (px3623), .I3 (px3439), .I4 (px3172)) ;
         defparam ix43824z28358.INIT = 32'h96696996;
    LUT6 ix43824z34719 (.O (px3035), .I0 (nx12903z176), .I1 (nx12903z180), .I2 (
         nx12903z174), .I3 (nx12903z178), .I4 (nx12903z182), .I5 (nx12903z172)
         ) ;
         defparam ix43824z34719.INIT = 64'hD11D3EA27CCB8274;
    (* HLUTNM = "LUT62_1_2" *)
    LUT5 ix35956z39819 (.O (px3036), .I0 (\plaintext(28)  ), .I1 (nx37232z9), .I2 (
         px3638), .I3 (px3442), .I4 (px3191)) ;
         defparam ix35956z39819.INIT = 32'h69969669;
    LUT6 ix12903z28592 (.O (nx12903z269), .I0 (\p_key_samp(6)  ), .I1 (
         nx12903z270), .I2 (nx15291z36), .I3 (nx13298z60), .I4 (nx12903z121), .I5 (
         nx12903z271)) ;
         defparam ix12903z28592.INIT = 64'h6996966996696996;
    LUT6 ix12903z48216 (.O (nx12903z271), .I0 (nx12903z272), .I1 (nx12903z273), 
         .I2 (nx12903z274), .I3 (nx12903z275), .I4 (nx12903z276), .I5 (
         nx12903z278)) ;
         defparam ix12903z48216.INIT = 64'hC3C4256B9C93B63C;
    (* HLUTNM = "LUT62_1_18" *)
    LUT5 ix43824z39822 (.O (nx43824z4), .I0 (\plaintext(52)  ), .I1 (nx36228z8)
         , .I2 (nx15291z36), .I3 (nx13298z60), .I4 (nx12903z121)) ;
         defparam ix43824z39822.INIT = 32'h69969669;
    LUT6 ix44815z28415 (.O (px3041), .I0 (nx12903z197), .I1 (nx12903z199), .I2 (
         nx12903z195), .I3 (nx12903z205), .I4 (nx12903z203), .I5 (nx12903z201)
         ) ;
         defparam ix44815z28415.INIT = 64'h6678B1CE798969D0;
    LUT6 ix12903z40013 (.O (nx12903z201), .I0 (\plaintext(31)  ), .I1 (
         \p_key_samp(62)  ), .I2 (nx28253z2), .I3 (px3562), .I4 (px3373), .I5 (
         px3112)) ;
         defparam ix12903z40013.INIT = 64'h9669699669969669;
    LUT6 ix12903z28540 (.O (nx12903z203), .I0 (\p_plaintext(39)  ), .I1 (
         \p_key_samp(29)  ), .I2 (px3781), .I3 (px3559), .I4 (px3353), .I5 (
         px3109)) ;
         defparam ix12903z28540.INIT = 64'h6996966996696996;
    LUT6 ix12903z28542 (.O (nx12903z205), .I0 (\plaintext(7)  ), .I1 (
         \p_key_samp(31)  ), .I2 (nx34235z6), .I3 (px3587), .I4 (px3304), .I5 (
         px3068)) ;
         defparam ix12903z28542.INIT = 64'h6996966996696996;
    LUT6 ix12903z28532 (.O (nx12903z195), .I0 (\plaintext(15)  ), .I1 (
         \p_key_samp(12)  ), .I2 (nx15291z18), .I3 (nx13298z54), .I4 (nx32966z9)
         , .I5 (nx12903z196)) ;
         defparam ix12903z28532.INIT = 64'h6996966996696996;
    LUT6 ix12903z27577 (.O (nx12903z196), .I0 (nx12903z100), .I1 (nx12903z103), 
         .I2 (nx12903z95), .I3 (nx12903z96), .I4 (nx12903z102), .I5 (nx12903z98)
         ) ;
         defparam ix12903z27577.INIT = 64'hC35AD2389C3565DA;
    (* HLUTNM = "LUT62_1_52" *)
    LUT4 ix43816z28368 (.O (nx43816z30), .I0 (\plaintext(15)  ), .I1 (nx15291z18
         ), .I2 (nx13298z54), .I3 (nx32966z9)) ;
         defparam ix43816z28368.INIT = 16'h6996;
    LUT6 ix12903z40011 (.O (nx12903z199), .I0 (\plaintext(23)  ), .I1 (
         \p_key_samp(22)  ), .I2 (nx15291z24), .I3 (nx13298z50), .I4 (nx32966z7)
         , .I5 (nx12903z200)) ;
         defparam ix12903z40011.INIT = 64'h9669699669969669;
    LUT6 ix12903z51289 (.O (nx12903z200), .I0 (nx12903z156), .I1 (nx12903z157), 
         .I2 (nx12903z158), .I3 (nx12903z159), .I4 (nx12903z161), .I5 (
         nx12903z162)) ;
         defparam ix12903z51289.INIT = 64'h7D6992C9B285C276;
    (* HLUTNM = "LUT62_1_53" *)
    LUT4 ix43816z39846 (.O (nx43816z33), .I0 (\plaintext(23)  ), .I1 (nx15291z24
         ), .I2 (nx13298z50), .I3 (nx32966z7)) ;
         defparam ix43816z39846.INIT = 16'h9669;
    LUT6 ix12903z28534 (.O (nx12903z197), .I0 (\plaintext(57)  ), .I1 (
         \p_key_samp(7)  ), .I2 (nx34235z21), .I3 (px3596), .I4 (px3307), .I5 (
         px3073)) ;
         defparam ix12903z28534.INIT = 64'h6996966996696996;
    (* HLUTNM = "LUT62_1_3" *)
    LUT5 ix37946z28344 (.O (px3052), .I0 (plaintext[4]), .I1 (nx36228z6), .I2 (
         px3626), .I3 (px3433), .I4 (px3183)) ;
         defparam ix37946z28344.INIT = 32'h96696996;
    LUT6 ix12903z21021 (.O (px3054), .I0 (nx12903z243), .I1 (nx12903z248), .I2 (
         nx12903z249), .I3 (nx12903z245), .I4 (nx12903z250), .I5 (nx12903z247)
         ) ;
         defparam ix12903z21021.INIT = 64'h96A999697C434BB4;
    (* HLUTNM = "LUT62_1_13" *)
    LUT5 ix43820z28347 (.O (nx43820z5), .I0 (\plaintext(36)  ), .I1 (nx37232z11)
         , .I2 (px3635), .I3 (px3436), .I4 (px3197)) ;
         defparam ix43820z28347.INIT = 32'h96696996;
    LUT6 ix42825z37099 (.O (px3057), .I0 (nx12903z340), .I1 (nx12903z345), .I2 (
         nx12903z342), .I3 (px3089), .I4 (px3076), .I5 (px3059)) ;
         defparam ix42825z37099.INIT = 64'h9E91661E960D8B75;
    LUT6 ix37952z61247 (.O (px3058), .I0 (nx12903z340), .I1 (nx12903z345), .I2 (
         nx12903z342), .I3 (px3089), .I4 (px3076), .I5 (px3059)) ;
         defparam ix37952z61247.INIT = 64'hCA3C75A230D6EA1D;
    LUT6 ix42825z38907 (.O (px3060), .I0 (nx12903z272), .I1 (nx12903z273), .I2 (
         nx12903z274), .I3 (nx12903z275), .I4 (nx12903z276), .I5 (nx12903z278)
         ) ;
         defparam ix42825z38907.INIT = 64'hB59C6CD24B599227;
    LUT6 ix12903z40076 (.O (nx12903z278), .I0 (\plaintext(41)  ), .I1 (
         \p_key_samp(2)  ), .I2 (nx34235z8), .I3 (nx13298z65), .I4 (nx12903z77)
         , .I5 (nx12903z279)) ;
         defparam ix12903z40076.INIT = 64'h9669699669969669;
    LUT6 ix12903z40065 (.O (nx12903z279), .I0 (nx12903z106), .I1 (nx12903z108), 
         .I2 (nx12903z110), .I3 (nx12903z112), .I4 (nx12903z113), .I5 (
         nx12903z114)) ;
         defparam ix12903z40065.INIT = 64'h66F91E41A156965D;
    (* HLUTNM = "LUT62_1_49" *)
    LUT4 ix42825z40005 (.O (nx42825z250), .I0 (\plaintext(41)  ), .I1 (nx34235z8
         ), .I2 (nx13298z65), .I3 (nx12903z77)) ;
         defparam ix42825z40005.INIT = 16'h9669;
    LUT6 ix12903z28599 (.O (nx12903z276), .I0 (\plaintext(49)  ), .I1 (
         \p_key_samp(51)  ), .I2 (nx34235z4), .I3 (nx13298z62), .I4 (nx12903z79)
         , .I5 (nx12903z277)) ;
         defparam ix12903z28599.INIT = 64'h6996966996696996;
    LUT6 ix12903z29437 (.O (nx12903z277), .I0 (nx12903z89), .I1 (nx12903z86), .I2 (
         nx12903z84), .I3 (nx12903z91), .I4 (nx12903z87), .I5 (nx12903z92)) ;
         defparam ix12903z29437.INIT = 64'h49DAB32986316CDB;
    (* HLUTNM = "LUT62_1_42" *)
    LUT4 ix42825z28527 (.O (nx42825z244), .I0 (\plaintext(49)  ), .I1 (nx34235z4
         ), .I2 (nx13298z62), .I3 (nx12903z79)) ;
         defparam ix42825z28527.INIT = 16'h6996;
    LUT6 ix12903z28598 (.O (nx12903z275), .I0 (\plaintext(7)  ), .I1 (
         \p_key_samp(19)  ), .I2 (nx34235z6), .I3 (px3587), .I4 (px3304), .I5 (
         px3068)) ;
         defparam ix12903z28598.INIT = 64'h6996966996696996;
    LUT6 ix12903z33949 (.O (px3068), .I0 (nx12903z117), .I1 (nx12903z118), .I2 (
         nx12903z119), .I3 (nx12903z120), .I4 (nx12903z122), .I5 (nx12903z124)
         ) ;
         defparam ix12903z33949.INIT = 64'hD487691E23C87EB4;
    (* HLUTNM = "LUT62_1_33" *)
    LUT4 ix38950z28344 (.O (px3069), .I0 (\plaintext(7)  ), .I1 (nx34235z6), .I2 (
         px3587), .I3 (px3304)) ;
         defparam ix38950z28344.INIT = 16'h6996;
    LUT6 ix12903z40072 (.O (nx12903z274), .I0 (\plaintext(25)  ), .I1 (
         \p_key_samp(33)  ), .I2 (nx34235z31), .I3 (px3590), .I4 (px3335), .I5 (
         px3151)) ;
         defparam ix12903z40072.INIT = 64'h9669699669969669;
    LUT6 ix12903z28596 (.O (nx12903z273), .I0 (\plaintext(33)  ), .I1 (
         \p_key_samp(1)  ), .I2 (nx34235z10), .I3 (px3584), .I4 (px3332), .I5 (
         px3154)) ;
         defparam ix12903z28596.INIT = 64'h6996966996696996;
    LUT6 ix12903z28595 (.O (nx12903z272), .I0 (\plaintext(57)  ), .I1 (
         \p_key_samp(58)  ), .I2 (nx34235z21), .I3 (px3596), .I4 (px3307), .I5 (
         px3073)) ;
         defparam ix12903z28595.INIT = 64'h6996966996696996;
    LUT6 ix12903z32645 (.O (px3073), .I0 (nx12903z142), .I1 (nx12903z143), .I2 (
         nx12903z144), .I3 (nx12903z146), .I4 (nx12903z148), .I5 (nx12903z149)
         ) ;
         defparam ix12903z32645.INIT = 64'hC93665C9B69479A4;
    (* HLUTNM = "LUT62_1_34" *)
    LUT4 ix39942z28344 (.O (px3074), .I0 (\plaintext(57)  ), .I1 (nx34235z21), .I2 (
         px3596), .I3 (px3307)) ;
         defparam ix39942z28344.INIT = 16'h6996;
    (* HLUTNM = "LUT62_1_8" *)
    LUT5 ix42825z28521 (.O (nx42825z238), .I0 (\plaintext(38)  ), .I1 (
         nx63157z36), .I2 (px3726), .I3 (px3582), .I4 (px3296)) ;
         defparam ix42825z28521.INIT = 32'h96696996;
    LUT6 ix42825z11154 (.O (px3077), .I0 (nx12903z229), .I1 (nx12903z230), .I2 (
         nx12903z231), .I3 (nx12903z233), .I4 (nx12903z234), .I5 (nx12903z236)
         ) ;
         defparam ix42825z11154.INIT = 64'h36CACA36F86525CA;
    LUT6 ix12903z28567 (.O (nx12903z236), .I0 (plaintext[5]), .I1 (
         \p_key_samp(49)  ), .I2 (nx27254z7), .I3 (px3543), .I4 (px3341), .I5 (
         px3138)) ;
         defparam ix12903z28567.INIT = 64'h6996966996696996;
    LUT6 ix12903z40039 (.O (nx12903z234), .I0 (\plaintext(51)  ), .I1 (
         \p_key_samp(25)  ), .I2 (nx25263z8), .I3 (nx24265z37), .I4 (nx12903z20)
         , .I5 (nx12903z235)) ;
         defparam ix12903z40039.INIT = 64'h9669699669969669;
    LUT6 ix12903z28785 (.O (nx12903z235), .I0 (nx12903z84), .I1 (nx12903z86), .I2 (
         nx12903z91), .I3 (nx12903z92), .I4 (nx12903z89), .I5 (nx12903z87)) ;
         defparam ix12903z28785.INIT = 64'hCABC636C17716992;
    (* HLUTNM = "LUT62_1_48" *)
    LUT4 ix42825z39993 (.O (nx42825z234), .I0 (\plaintext(51)  ), .I1 (nx25263z8
         ), .I2 (nx24265z37), .I3 (nx12903z20)) ;
         defparam ix42825z39993.INIT = 16'h9669;
    LUT6 ix12903z28563 (.O (nx12903z233), .I0 (\plaintext(27)  ), .I1 (
         \p_key_samp(3)  ), .I2 (nx36228z2), .I3 (px3615), .I4 (px3425), .I5 (
         px3170)) ;
         defparam ix12903z28563.INIT = 64'h6996966996696996;
    LUT6 ix12903z28561 (.O (nx12903z231), .I0 (\plaintext(43)  ), .I1 (
         \p_key_samp(10)  ), .I2 (nx25263z6), .I3 (nx24265z26), .I4 (nx12903z22)
         , .I5 (nx12903z232)) ;
         defparam ix12903z28561.INIT = 64'h6996966996696996;
    LUT6 ix12903z9437 (.O (nx12903z232), .I0 (nx12903z143), .I1 (nx12903z144), .I2 (
         nx12903z146), .I3 (nx12903z148), .I4 (nx12903z149), .I5 (nx12903z142)
         ) ;
         defparam ix12903z9437.INIT = 64'hEC78C38D23961EE1;
    (* HLUTNM = "LUT62_1_41" *)
    LUT4 ix42825z28515 (.O (nx42825z230), .I0 (\plaintext(43)  ), .I1 (nx25263z6
         ), .I2 (nx24265z26), .I3 (nx12903z22)) ;
         defparam ix42825z28515.INIT = 16'h6996;
    LUT6 ix12903z28560 (.O (nx12903z230), .I0 (\plaintext(59)  ), .I1 (
         \p_key_samp(27)  ), .I2 (nx27254z4), .I3 (px3546), .I4 (px3338), .I5 (
         px3160)) ;
         defparam ix12903z28560.INIT = 64'h6996966996696996;
    LUT6 ix12903z40034 (.O (nx12903z229), .I0 (\plaintext(35)  ), .I1 (
         \p_key_samp(52)  ), .I2 (nx39226z2), .I3 (px3652), .I4 (px3408), .I5 (
         px3245)) ;
         defparam ix12903z40034.INIT = 64'h9669699669969669;
    (* HLUTNM = "LUT62_1_7" *)
    LUT5 ix42825z28509 (.O (nx42825z222), .I0 (\plaintext(30)  ), .I1 (
         nx63157z44), .I2 (px3752), .I3 (px3523), .I4 (px3283)) ;
         defparam ix42825z28509.INIT = 32'h96696996;
    LUT6 ix61487z53854 (.O (px3090), .I0 (nx12903z357), .I1 (nx12903z359), .I2 (
         nx12903z362), .I3 (nx12903z361), .I4 (nx12903z358), .I5 (nx12903z364)
         ) ;
         defparam ix61487z53854.INIT = 64'h364E78A1D0E9CD36;
    LUT6 ix12903z28668 (.O (nx12903z364), .I0 (\p_plaintext(37)  ), .I1 (
         \p_key_samp(45)  ), .I2 (px3745), .I3 (px3514), .I4 (px3315), .I5 (
         px3092)) ;
         defparam ix12903z28668.INIT = 64'h6996966996696996;
    LUT6 ix12903z30802 (.O (px3092), .I0 (nx12903z95), .I1 (nx12903z96), .I2 (
         nx12903z98), .I3 (nx12903z100), .I4 (nx12903z102), .I5 (nx12903z103)) ;
         defparam ix12903z30802.INIT = 64'h56B8876969C3729C;
    (* HLUTNM = "LUT62_1_35" *)
    LUT4 ix41935z28344 (.O (px3093), .I0 (\p_plaintext(37)  ), .I1 (px3745), .I2 (
         px3514), .I3 (px3315)) ;
         defparam ix41935z28344.INIT = 16'h6996;
    LUT6 ix12903z28662 (.O (nx12903z358), .I0 (\plaintext(29)  ), .I1 (
         \p_key_samp(23)  ), .I2 (nx23267z2), .I3 (px3511), .I4 (px3321), .I5 (
         px3095)) ;
         defparam ix12903z28662.INIT = 64'h6996966996696996;
    LUT6 ix12903z27508 (.O (px3095), .I0 (nx12903z142), .I1 (nx12903z143), .I2 (
         nx12903z144), .I3 (nx12903z146), .I4 (nx12903z148), .I5 (nx12903z149)
         ) ;
         defparam ix12903z27508.INIT = 64'h6E38396C9C6665C9;
    (* HLUTNM = "LUT62_1_36" *)
    LUT4 ix41938z28344 (.O (px3096), .I0 (\plaintext(29)  ), .I1 (nx23267z2), .I2 (
         px3511), .I3 (px3321)) ;
         defparam ix41938z28344.INIT = 16'h6996;
    LUT6 ix12903z28665 (.O (nx12903z361), .I0 (\plaintext(61)  ), .I1 (
         \p_key_samp(28)  ), .I2 (nx37232z2), .I3 (px3632), .I4 (px3392), .I5 (
         px3187)) ;
         defparam ix12903z28665.INIT = 64'h6996966996696996;
    LUT6 ix12903z28666 (.O (nx12903z362), .I0 (\plaintext(45)  ), .I1 (
         \p_key_samp(46)  ), .I2 (nx16289z7), .I3 (nx7312z12), .I4 (nx12903z36)
         , .I5 (nx12903z363)) ;
         defparam ix12903z28666.INIT = 64'h6996966996696996;
    LUT6 ix12903z40910 (.O (nx12903z363), .I0 (nx12903z159), .I1 (nx12903z158), 
         .I2 (nx12903z161), .I3 (nx12903z162), .I4 (nx12903z157), .I5 (
         nx12903z156)) ;
         defparam ix12903z40910.INIT = 64'hE44B279663B49969;
    (* HLUTNM = "LUT62_1_47" *)
    LUT4 ix42825z39975 (.O (nx42825z207), .I0 (\plaintext(45)  ), .I1 (nx16289z7
         ), .I2 (nx7312z12), .I3 (nx12903z36)) ;
         defparam ix42825z39975.INIT = 16'h9669;
    LUT6 ix12903z28663 (.O (nx12903z359), .I0 (\plaintext(53)  ), .I1 (
         \p_key_samp(55)  ), .I2 (nx16289z10), .I3 (nx7312z17), .I4 (nx12903z31)
         , .I5 (nx12903z360)) ;
         defparam ix12903z28663.INIT = 64'h6996966996696996;
    LUT6 ix12903z37083 (.O (nx12903z360), .I0 (nx12903z16), .I1 (nx12903z26), .I2 (
         nx12903z28), .I3 (nx12903z38), .I4 (nx12903z48), .I5 (nx12903z50)) ;
         defparam ix12903z37083.INIT = 64'hB99655A699438A79;
    (* HLUTNM = "LUT62_1_46" *)
    LUT4 ix42825z39972 (.O (nx42825z203), .I0 (\plaintext(53)  ), .I1 (
         nx16289z10), .I2 (nx7312z17), .I3 (nx12903z31)) ;
         defparam ix42825z39972.INIT = 16'h9669;
    LUT6 ix12903z40136 (.O (nx12903z357), .I0 (plaintext[3]), .I1 (
         \p_key_samp(5)  ), .I2 (nx38222z2), .I3 (px3649), .I4 (px3405), .I5 (
         px3221)) ;
         defparam ix12903z40136.INIT = 64'h9669699669969669;
    (* HLUTNM = "LUT62_1_6" *)
    LUT5 ix42825z28493 (.O (nx42825z198), .I0 (plaintext[0]), .I1 (nx63157z28), 
         .I2 (px3739), .I3 (px3506), .I4 (px3313)) ;
         defparam ix42825z28493.INIT = 32'h96696996;
    LUT6 ix12903z28647 (.O (nx12903z342), .I0 (\p_key_samp(28)  ), .I1 (
         nx12903z343), .I2 (nx37234z7), .I3 (nx11304z6), .I4 (nx12903z88), .I5 (
         nx12903z344)) ;
         defparam ix12903z28647.INIT = 64'h6996966996696996;
    LUT6 ix12903z27771 (.O (nx12903z344), .I0 (nx12903z243), .I1 (nx12903z248), 
         .I2 (nx12903z249), .I3 (nx12903z245), .I4 (nx12903z250), .I5 (
         nx12903z247)) ;
         defparam ix12903z27771.INIT = 64'h87D179C7D12E6628;
    LUT6 ix12903z28575 (.O (nx12903z247), .I0 (\p_plaintext(39)  ), .I1 (
         \p_key_samp(54)  ), .I2 (px3781), .I3 (px3559), .I4 (px3353), .I5 (
         px3109)) ;
         defparam ix12903z28575.INIT = 64'h6996966996696996;
    LUT6 ix12903z28111 (.O (px3109), .I0 (nx12903z16), .I1 (nx12903z26), .I2 (
         nx12903z28), .I3 (nx12903z38), .I4 (nx12903z48), .I5 (nx12903z50)) ;
         defparam ix12903z28111.INIT = 64'h21D99C47DA2967E8;
    (* HLUTNM = "LUT62_1_54" *)
    LUT4 ix44925z28344 (.O (px3110), .I0 (\p_plaintext(39)  ), .I1 (px3781), .I2 (
         px3559), .I3 (px3353)) ;
         defparam ix44925z28344.INIT = 16'h6996;
    LUT6 ix12903z40053 (.O (nx12903z250), .I0 (\plaintext(31)  ), .I1 (
         \p_key_samp(13)  ), .I2 (nx28253z2), .I3 (px3562), .I4 (px3373), .I5 (
         px3112)) ;
         defparam ix12903z40053.INIT = 64'h9669699669969669;
    LUT6 ix12903z55314 (.O (px3112), .I0 (nx12903z70), .I1 (nx12903z64), .I2 (
         nx12903z66), .I3 (nx12903z62), .I4 (nx12903z68), .I5 (nx12903z80)) ;
         defparam ix12903z55314.INIT = 64'hE92E25D223E9D22D;
    (* HLUTNM = "LUT62_1_55" *)
    LUT4 ix44928z39819 (.O (px3113), .I0 (\plaintext(31)  ), .I1 (nx28253z2), .I2 (
         px3562), .I3 (px3373)) ;
         defparam ix44928z39819.INIT = 16'h9669;
    LUT6 ix12903z28573 (.O (nx12903z245), .I0 (\plaintext(47)  ), .I1 (
         \p_key_samp(15)  ), .I2 (nx15291z12), .I3 (nx13298z46), .I4 (nx12903z46
         ), .I5 (nx12903z246)) ;
         defparam ix12903z28573.INIT = 64'h6996966996696996;
    LUT6 ix12903z40772 (.O (nx12903z246), .I0 (nx12903z106), .I1 (nx12903z108), 
         .I2 (nx12903z110), .I3 (nx12903z112), .I4 (nx12903z113), .I5 (
         nx12903z114)) ;
         defparam ix12903z40772.INIT = 64'h94F26A9566C3993C;
    (* HLUTNM = "LUT62_1_39" *)
    LUT4 ix42825z28453 (.O (nx42825z140), .I0 (\plaintext(47)  ), .I1 (
         nx15291z12), .I2 (nx13298z46), .I3 (nx12903z46)) ;
         defparam ix42825z28453.INIT = 16'h6996;
    LUT6 ix12903z28577 (.O (nx12903z249), .I0 (p_nbus_plaintext[63]), .I1 (
         \p_key_samp(4)  ), .I2 (nx63157z2), .I3 (px3724), .I4 (px3504), .I5 (
         px3281)) ;
         defparam ix12903z28577.INIT = 64'h6996966996696996;
    LUT6 ix12903z40051 (.O (nx12903z248), .I0 (\p_plaintext(63)  ), .I1 (
         \p_key_samp(63)  ), .I2 (nx29253z2), .I3 (px3565), .I4 (px3359), .I5 (
         px3119)) ;
         defparam ix12903z40051.INIT = 64'h9669699669969669;
    LUT6 ix12903z39556 (.O (px3119), .I0 (nx12903z156), .I1 (nx12903z157), .I2 (
         nx12903z158), .I3 (nx12903z159), .I4 (nx12903z161), .I5 (nx12903z162)
         ) ;
         defparam ix12903z39556.INIT = 64'h54B2A36D79C394CA;
    (* HLUTNM = "LUT62_1_56" *)
    LUT4 ix45922z39819 (.O (px3120), .I0 (\p_plaintext(63)  ), .I1 (nx29253z2), 
         .I2 (px3565), .I3 (px3359)) ;
         defparam ix45922z39819.INIT = 16'h9669;
    LUT6 ix12903z28571 (.O (nx12903z243), .I0 (\plaintext(55)  ), .I1 (
         \p_key_samp(37)  ), .I2 (nx15291z8), .I3 (nx13298z39), .I4 (nx12903z41)
         , .I5 (nx12903z244)) ;
         defparam ix12903z28571.INIT = 64'h6996966996696996;
    LUT6 ix12903z17056 (.O (nx12903z244), .I0 (nx12903z142), .I1 (nx12903z143), 
         .I2 (nx12903z144), .I3 (nx12903z146), .I4 (nx12903z148), .I5 (
         nx12903z149)) ;
         defparam ix12903z17056.INIT = 64'h389EC36586793C9A;
    LUT6 ix12903z39965 (.O (nx12903z149), .I0 (\plaintext(58)  ), .I1 (
         \p_key_samp(9)  ), .I2 (nx34235z18), .I3 (px3705), .I4 (px3460), .I5 (
         px3232)) ;
         defparam ix12903z39965.INIT = 64'h9669699669969669;
    LUT6 ix12903z28489 (.O (nx12903z148), .I0 (\plaintext(32)  ), .I1 (
         \p_key_samp(18)  ), .I2 (nx39226z15), .I3 (px3665), .I4 (px3421), .I5 (
         px3278)) ;
         defparam ix12903z28489.INIT = 64'h6996966996696996;
    LUT6 ix12903z28487 (.O (nx12903z146), .I0 (\plaintext(8)  ), .I1 (
         \p_key_samp(36)  ), .I2 (nx34235z25), .I3 (nx24265z31), .I4 (nx337z6), 
         .I5 (nx12903z147)) ;
         defparam ix12903z28487.INIT = 64'h6996966996696996;
    LUT6 ix12903z41194 (.O (nx12903z147), .I0 (nx12903z30), .I1 (nx12903z32), .I2 (
         nx12903z33), .I3 (nx12903z34), .I4 (nx12903z35), .I5 (nx12903z37)) ;
         defparam ix12903z41194.INIT = 64'hED16146658E79B38;
    (* HLUTNM = "LUT62_1_38" *)
    LUT4 ix42825z28425 (.O (nx42825z100), .I0 (\plaintext(8)  ), .I1 (nx34235z25
         ), .I2 (nx24265z31), .I3 (nx337z6)) ;
         defparam ix42825z28425.INIT = 16'h6996;
    LUT6 ix12903z28485 (.O (nx12903z144), .I0 (\plaintext(16)  ), .I1 (
         \p_key_samp(42)  ), .I2 (nx34235z28), .I3 (nx24265z33), .I4 (nx337z4), 
         .I5 (nx12903z145)) ;
         defparam ix12903z28485.INIT = 64'h6996966996696996;
    LUT6 ix12903z40951 (.O (nx12903z145), .I0 (nx12903z72), .I1 (nx12903z73), .I2 (
         nx12903z74), .I3 (nx12903z75), .I4 (nx12903z76), .I5 (nx12903z78)) ;
         defparam ix12903z40951.INIT = 64'h51ADE51A2EE19A47;
    (* HLUTNM = "LUT62_1_29" *)
    LUT4 ix42825z39915 (.O (nx42825z120), .I0 (\plaintext(16)  ), .I1 (
         nx34235z28), .I2 (nx24265z33), .I3 (nx337z4)) ;
         defparam ix42825z39915.INIT = 16'h9669;
    LUT6 ix12903z28484 (.O (nx12903z143), .I0 (\plaintext(24)  ), .I1 (
         \p_key_samp(27)  ), .I2 (nx39226z17), .I3 (px3657), .I4 (px3410), .I5 (
         px3261)) ;
         defparam ix12903z28484.INIT = 64'h6996966996696996;
    LUT6 ix12903z28623 (.O (nx12903z142), .I0 (plaintext[6]), .I1 (
         \p_key_samp(49)  ), .I2 (nx44209z2), .I3 (px3702), .I4 (px3451), .I5 (
         px3235)) ;
         defparam ix12903z28623.INIT = 64'h6996966996696996;
    (* HLUTNM = "LUT62_1_44" *)
    LUT4 ix42825z39897 (.O (nx42825z97), .I0 (\plaintext(55)  ), .I1 (nx15291z8)
         , .I2 (nx13298z39), .I3 (nx12903z41)) ;
         defparam ix42825z39897.INIT = 16'h9669;
    (* HLUTNM = "LUT62_1_9" *)
    LUT5 ix42825z39894 (.O (nx42825z94), .I0 (\plaintext(14)  ), .I1 (nx63157z12
         ), .I2 (nx37234z7), .I3 (nx11304z6), .I4 (nx12903z88)) ;
         defparam ix42825z39894.INIT = 32'h69969669;
    LUT6 ix12903z28650 (.O (nx12903z345), .I0 (\p_key_samp(23)  ), .I1 (
         nx12903z296), .I2 (nx27254z2), .I3 (px3536), .I4 (px3330), .I5 (px3136)
         ) ;
         defparam ix12903z28650.INIT = 64'h6996966996696996;
    LUT6 ix12903z41218 (.O (px3136), .I0 (nx12903z176), .I1 (nx12903z180), .I2 (
         nx12903z174), .I3 (nx12903z178), .I4 (nx12903z182), .I5 (nx12903z172)
         ) ;
         defparam ix12903z41218.INIT = 64'hB84BC3A865B69AD1;
    LUT6 ix12903z28511 (.O (nx12903z172), .I0 (plaintext[5]), .I1 (
         \p_key_samp(57)  ), .I2 (nx27254z7), .I3 (px3543), .I4 (px3341), .I5 (
         px3138)) ;
         defparam ix12903z28511.INIT = 64'h6996966996696996;
    LUT6 ix12903z14568 (.O (px3138), .I0 (nx12903z156), .I1 (nx12903z157), .I2 (
         nx12903z158), .I3 (nx12903z159), .I4 (nx12903z161), .I5 (nx12903z162)
         ) ;
         defparam ix12903z14568.INIT = 64'hB65BC8E42CD1331E;
    LUT6 ix12903z39978 (.O (nx12903z162), .I0 (\plaintext(18)  ), .I1 (
         \p_key_samp(51)  ), .I2 (nx29253z8), .I3 (nx24265z20), .I4 (nx4319z5), 
         .I5 (nx12903z163)) ;
         defparam ix12903z39978.INIT = 64'h9669699669969669;
    LUT6 ix12903z41435 (.O (nx12903z163), .I0 (nx12903z21), .I1 (nx12903z23), .I2 (
         nx12903z25), .I3 (nx12903z24), .I4 (nx12903z18), .I5 (nx12903z19)) ;
         defparam ix12903z41435.INIT = 64'hE40F935A63F49C19;
    (* HLUTNM = "LUT62_1_21" *)
    LUT4 ix42825z39978 (.O (nx42825z210), .I0 (\plaintext(18)  ), .I1 (nx29253z8
         ), .I2 (nx24265z20), .I3 (nx4319z5)) ;
         defparam ix42825z39978.INIT = 16'h9669;
    LUT6 ix12903z28502 (.O (nx12903z161), .I0 (plaintext[4]), .I1 (
         \p_key_samp(10)  ), .I2 (nx36228z6), .I3 (px3626), .I4 (px3433), .I5 (
         px3183)) ;
         defparam ix12903z28502.INIT = 64'h6996966996696996;
    LUT6 ix12903z39975 (.O (nx12903z159), .I0 (\plaintext(10)  ), .I1 (
         \p_key_samp(3)  ), .I2 (nx29253z10), .I3 (nx24265z23), .I4 (nx4319z3), 
         .I5 (nx12903z160)) ;
         defparam ix12903z39975.INIT = 64'h9669699669969669;
    LUT6 ix12903z38191 (.O (nx12903z160), .I0 (nx12903z45), .I1 (nx12903z44), .I2 (
         nx12903z42), .I3 (nx12903z40), .I4 (nx12903z43), .I5 (nx12903z47)) ;
         defparam ix12903z38191.INIT = 64'hD919A16D21EE8F70;
    (* HLUTNM = "LUT62_1_22" *)
    LUT4 ix42825z39981 (.O (nx42825z217), .I0 (\plaintext(10)  ), .I1 (
         nx29253z10), .I2 (nx24265z23), .I3 (nx4319z3)) ;
         defparam ix42825z39981.INIT = 16'h9669;
    LUT6 ix12903z28499 (.O (nx12903z158), .I0 (\plaintext(26)  ), .I1 (
         \p_key_samp(33)  ), .I2 (nx45210z2), .I3 (px3716), .I4 (px3454), .I5 (
         px3226)) ;
         defparam ix12903z28499.INIT = 64'h6996966996696996;
    LUT6 ix12903z28498 (.O (nx12903z157), .I0 (\plaintext(60)  ), .I1 (
         \p_key_samp(52)  ), .I2 (nx36228z10), .I3 (px3623), .I4 (px3439), .I5 (
         px3172)) ;
         defparam ix12903z28498.INIT = 64'h6996966996696996;
    LUT6 ix12903z39972 (.O (nx12903z156), .I0 (\plaintext(34)  ), .I1 (
         \p_key_samp(34)  ), .I2 (nx41222z2), .I3 (px3688), .I4 (px3448), .I5 (
         px3229)) ;
         defparam ix12903z39972.INIT = 64'h9669699669969669;
    (* HLUTNM = "LUT62_1_57" *)
    LUT4 ix47925z28344 (.O (px3149), .I0 (plaintext[5]), .I1 (nx27254z7), .I2 (
         px3543), .I3 (px3341)) ;
         defparam ix47925z28344.INIT = 16'h6996;
    LUT6 ix12903z39996 (.O (nx12903z182), .I0 (\plaintext(25)  ), .I1 (
         \p_key_samp(35)  ), .I2 (nx34235z31), .I3 (px3590), .I4 (px3335), .I5 (
         px3151)) ;
         defparam ix12903z39996.INIT = 64'h9669699669969669;
    LUT6 ix12903z39322 (.O (px3151), .I0 (nx12903z95), .I1 (nx12903z96), .I2 (
         nx12903z98), .I3 (nx12903z100), .I4 (nx12903z102), .I5 (nx12903z103)) ;
         defparam ix12903z39322.INIT = 64'hC5363AC964B993C6;
    (* HLUTNM = "LUT62_1_58" *)
    LUT4 ix48915z28344 (.O (px3152), .I0 (\plaintext(25)  ), .I1 (nx34235z31), .I2 (
         px3590), .I3 (px3335)) ;
         defparam ix48915z28344.INIT = 16'h6996;
    LUT6 ix12903z28517 (.O (nx12903z178), .I0 (\plaintext(33)  ), .I1 (
         \p_key_samp(26)  ), .I2 (nx34235z10), .I3 (px3584), .I4 (px3332), .I5 (
         px3154)) ;
         defparam ix12903z28517.INIT = 64'h6996966996696996;
    LUT6 ix12903z12710 (.O (px3154), .I0 (nx12903z62), .I1 (nx12903z64), .I2 (
         nx12903z80), .I3 (nx12903z70), .I4 (nx12903z66), .I5 (nx12903z68)) ;
         defparam ix12903z12710.INIT = 64'hC39A34697C232BD6;
    (* HLUTNM = "LUT62_1_59" *)
    LUT4 ix48918z28344 (.O (px3155), .I0 (\plaintext(33)  ), .I1 (nx34235z10), .I2 (
         px3584), .I3 (px3332)) ;
         defparam ix48918z28344.INIT = 16'h6996;
    LUT6 ix12903z28513 (.O (nx12903z174), .I0 (\plaintext(9)  ), .I1 (
         \p_key_samp(44)  ), .I2 (nx27254z9), .I3 (nx13298z5), .I4 (nx35956z4), 
         .I5 (nx12903z175)) ;
         defparam ix12903z28513.INIT = 64'h6996966996696996;
    LUT6 ix12903z47706 (.O (nx12903z175), .I0 (nx12903z117), .I1 (nx12903z118), 
         .I2 (nx12903z119), .I3 (nx12903z120), .I4 (nx12903z122), .I5 (
         nx12903z124)) ;
         defparam ix12903z47706.INIT = 64'h87DB4C31D269B48E;
    (* HLUTNM = "LUT62_1_40" *)
    LUT4 ix42825z28475 (.O (nx42825z168), .I0 (\plaintext(9)  ), .I1 (nx27254z9)
         , .I2 (nx13298z5), .I3 (nx35956z4)) ;
         defparam ix42825z28475.INIT = 16'h6996;
    LUT6 ix12903z28519 (.O (nx12903z180), .I0 (\plaintext(59)  ), .I1 (
         \p_key_samp(17)  ), .I2 (nx27254z4), .I3 (px3546), .I4 (px3338), .I5 (
         px3160)) ;
         defparam ix12903z28519.INIT = 64'h6996966996696996;
    LUT6 ix12903z52268 (.O (px3160), .I0 (nx12903z113), .I1 (nx12903z108), .I2 (
         nx12903z106), .I3 (nx12903z114), .I4 (nx12903z110), .I5 (nx12903z112)
         ) ;
         defparam ix12903z52268.INIT = 64'hC2793DA239C6C65A;
    (* HLUTNM = "LUT62_1_60" *)
    LUT4 ix49911z39819 (.O (px3161), .I0 (\plaintext(59)  ), .I1 (nx27254z4), .I2 (
         px3546), .I3 (px3338)) ;
         defparam ix49911z39819.INIT = 16'h9669;
    LUT6 ix12903z28515 (.O (nx12903z176), .I0 (\plaintext(17)  ), .I1 (
         \p_key_samp(50)  ), .I2 (nx27254z11), .I3 (nx13298z9), .I4 (nx35956z6)
         , .I5 (nx12903z177)) ;
         defparam ix12903z28515.INIT = 64'h6996966996696996;
    LUT6 ix12903z59187 (.O (nx12903z177), .I0 (nx12903z16), .I1 (nx12903z26), .I2 (
         nx12903z28), .I3 (nx12903z38), .I4 (nx12903z48), .I5 (nx12903z50)) ;
         defparam ix12903z59187.INIT = 64'h69614B9E3C6AE165;
    (* HLUTNM = "LUT62_1_45" *)
    LUT4 ix42825z39959 (.O (nx42825z183), .I0 (\plaintext(17)  ), .I1 (
         nx27254z11), .I2 (nx13298z9), .I3 (nx35956z6)) ;
         defparam ix42825z39959.INIT = 16'h9669;
    (* HLUTNM = "LUT62_1_5" *)
    LUT5 ix42825z28470 (.O (nx42825z163), .I0 (\plaintext(56)  ), .I1 (
         nx63157z20), .I2 (nx27254z2), .I3 (px3536), .I4 (px3330)) ;
         defparam ix42825z28470.INIT = 32'h96696996;
    LUT6 ix12903z28645 (.O (nx12903z340), .I0 (\p_key_samp(38)  ), .I1 (
         nx12903z341), .I2 (nx37234z3), .I3 (nx11304z3), .I4 (nx12903z4), .I5 (
         nx12903z13)) ;
         defparam ix12903z28645.INIT = 64'h6996966996696996;
    (* HLUTNM = "LUT62_1_4" *)
    LUT5 ix42825z28347 (.O (nx42825z4), .I0 (\plaintext(22)  ), .I1 (nx63157z4)
         , .I2 (nx37234z3), .I3 (nx11304z3), .I4 (nx12903z4)) ;
         defparam ix42825z28347.INIT = 32'h96696996;
    LUT6 ix12903z29337 (.O (nx12903z13), .I0 (nx12903z14), .I1 (nx12903z60), .I2 (
         nx12903z82), .I3 (nx12903z93), .I4 (nx12903z104), .I5 (nx12903z115)) ;
         defparam ix12903z29337.INIT = 64'h65A63099F21C6D6B;
    LUT6 ix12903z28458 (.O (nx12903z115), .I0 (\plaintext(27)  ), .I1 (
         \p_key_samp(41)  ), .I2 (nx36228z2), .I3 (px3615), .I4 (px3425), .I5 (
         px3170)) ;
         defparam ix12903z28458.INIT = 64'h6996966996696996;
    LUT6 ix12903z12973 (.O (px3170), .I0 (nx12903z117), .I1 (nx12903z118), .I2 (
         nx12903z119), .I3 (nx12903z120), .I4 (nx12903z122), .I5 (nx12903z124)
         ) ;
         defparam ix12903z12973.INIT = 64'h1EB2D967B4C32D18;
    LUT6 ix12903z28467 (.O (nx12903z124), .I0 (\plaintext(60)  ), .I1 (
         \p_key_samp(20)  ), .I2 (nx36228z10), .I3 (px3623), .I4 (px3439), .I5 (
         px3172)) ;
         defparam ix12903z28467.INIT = 64'h6996966996696996;
    LUT6 ix12903z61108 (.O (px3172), .I0 (nx12903z52), .I1 (nx12903z53), .I2 (
         nx12903z54), .I3 (nx12903z56), .I4 (nx12903z57), .I5 (nx12903z59)) ;
         defparam ix12903z61108.INIT = 64'h5B2626D949D6E916;
    (* HLUTNM = "LUT62_1_17" *)
    LUT4 ix50910z39819 (.O (px3173), .I0 (\plaintext(60)  ), .I1 (nx36228z10), .I2 (
         px3623), .I3 (px3439)) ;
         defparam ix50910z39819.INIT = 16'h9669;
    LUT6 ix12903z28465 (.O (nx12903z122), .I0 (\plaintext(44)  ), .I1 (
         \p_key_samp(38)  ), .I2 (nx36228z4), .I3 (nx15291z38), .I4 (nx13298z70)
         , .I5 (nx12903z123)) ;
         defparam ix12903z28465.INIT = 64'h6996966996696996;
    LUT6 ix12903z59608 (.O (nx12903z123), .I0 (nx12903z7), .I1 (nx12903z5), .I2 (
         nx12903z10), .I3 (nx12903z9), .I4 (nx12903z11), .I5 (nx12903z12)) ;
         defparam ix12903z59608.INIT = 64'h8DB65A619649E33C;
    (* HLUTNM = "LUT62_1_16" *)
    LUT4 ix42825z39953 (.O (nx42825z173), .I0 (\plaintext(44)  ), .I1 (nx36228z4
         ), .I2 (nx15291z38), .I3 (nx13298z70)) ;
         defparam ix42825z39953.INIT = 16'h9669;
    LUT6 ix12903z39938 (.O (nx12903z120), .I0 (\plaintext(52)  ), .I1 (
         \p_key_samp(47)  ), .I2 (nx36228z8), .I3 (nx15291z36), .I4 (nx13298z60)
         , .I5 (nx12903z121)) ;
         defparam ix12903z39938.INIT = 64'h9669699669969669;
    LUT6 ix12903z28659 (.O (nx12903z121), .I0 (nx12903z72), .I1 (nx12903z73), .I2 (
         nx12903z74), .I3 (nx12903z75), .I4 (nx12903z76), .I5 (nx12903z78)) ;
         defparam ix12903z28659.INIT = 64'h34976D6699A86A59;
    (* HLUTNM = "LUT62_1_18" *)
    LUT4 ix42825z39956 (.O (nx42825z177), .I0 (\plaintext(52)  ), .I1 (nx36228z8
         ), .I2 (nx15291z36), .I3 (nx13298z60)) ;
         defparam ix42825z39956.INIT = 16'h9669;
    LUT6 ix12903z39937 (.O (nx12903z119), .I0 (\plaintext(28)  ), .I1 (
         \p_key_samp(15)  ), .I2 (nx37232z9), .I3 (px3638), .I4 (px3442), .I5 (
         px3191)) ;
         defparam ix12903z39937.INIT = 64'h9669699669969669;
    LUT6 ix12903z28461 (.O (nx12903z118), .I0 (\plaintext(36)  ), .I1 (
         \p_key_samp(37)  ), .I2 (nx37232z11), .I3 (px3635), .I4 (px3436), .I5 (
         px3197)) ;
         defparam ix12903z28461.INIT = 64'h6996966996696996;
    LUT6 ix12903z28460 (.O (nx12903z117), .I0 (plaintext[4]), .I1 (
         \p_key_samp(62)  ), .I2 (nx36228z6), .I3 (px3626), .I4 (px3433), .I5 (
         px3183)) ;
         defparam ix12903z28460.INIT = 64'h6996966996696996;
    LUT6 ix37946z19163 (.O (px3183), .I0 (nx32966z3), .I1 (nx32966z4), .I2 (
         nx32966z5), .I3 (nx32966z6), .I4 (nx32966z8), .I5 (nx32966z10)) ;
         defparam ix37946z19163.INIT = 64'h35DE6942DE2645B8;
    (* HLUTNM = "LUT62_1_3" *)
    LUT4 ix51908z28344 (.O (px3184), .I0 (plaintext[4]), .I1 (nx36228z6), .I2 (
         px3626), .I3 (px3433)) ;
         defparam ix51908z28344.INIT = 16'h6996;
    (* HLUTNM = "LUT62_1_61" *)
    LUT4 ix51909z28344 (.O (px3185), .I0 (\plaintext(27)  ), .I1 (nx36228z2), .I2 (
         px3615), .I3 (px3425)) ;
         defparam ix51909z28344.INIT = 16'h6996;
    LUT6 ix12903z28447 (.O (nx12903z104), .I0 (\plaintext(61)  ), .I1 (
         \p_key_samp(60)  ), .I2 (nx37232z2), .I3 (px3632), .I4 (px3392), .I5 (
         px3187)) ;
         defparam ix12903z28447.INIT = 64'h6996966996696996;
    LUT6 ix12903z51424 (.O (px3187), .I0 (nx12903z106), .I1 (nx12903z108), .I2 (
         nx12903z110), .I3 (nx12903z112), .I4 (nx12903z113), .I5 (nx12903z114)
         ) ;
         defparam ix12903z51424.INIT = 64'hD3661CA9ACB1C356;
    LUT6 ix12903z39932 (.O (nx12903z114), .I0 (\plaintext(62)  ), .I1 (
         \p_key_samp(6)  ), .I2 (nx37232z13), .I3 (nx36230z11), .I4 (nx9305z10)
         , .I5 (px3216)) ;
         defparam ix12903z39932.INIT = 64'h9669699669969669;
    LUT6 ix12903z39931 (.O (nx12903z113), .I0 (plaintext[2]), .I1 (
         \p_key_samp(39)  ), .I2 (nx40221z2), .I3 (px3674), .I4 (px3483), .I5 (
         px3206)) ;
         defparam ix12903z39931.INIT = 64'h9669699669969669;
    LUT6 ix12903z39930 (.O (nx12903z112), .I0 (\plaintext(28)  ), .I1 (
         \p_key_samp(30)  ), .I2 (nx37232z9), .I3 (px3638), .I4 (px3442), .I5 (
         px3191)) ;
         defparam ix12903z39930.INIT = 64'h9669699669969669;
    LUT6 ix35956z16207 (.O (px3191), .I0 (nx35956z3), .I1 (nx35956z5), .I2 (
         nx35956z7), .I3 (nx35956z8), .I4 (nx35956z9), .I5 (nx35956z10)) ;
         defparam ix35956z16207.INIT = 64'hCAADB152C55B3A2C;
    (* HLUTNM = "LUT62_1_2" *)
    LUT4 ix52903z39819 (.O (px3192), .I0 (\plaintext(28)  ), .I1 (nx37232z9), .I2 (
         px3638), .I3 (px3442)) ;
         defparam ix52903z39819.INIT = 16'h9669;
    LUT6 ix12903z28453 (.O (nx12903z110), .I0 (\plaintext(20)  ), .I1 (
         \p_key_samp(13)  ), .I2 (nx37232z6), .I3 (nx36230z5), .I4 (nx9305z5), .I5 (
         nx12903z111)) ;
         defparam ix12903z28453.INIT = 64'h6996966996696996;
    LUT6 ix12903z55292 (.O (nx12903z111), .I0 (nx12903z18), .I1 (nx12903z21), .I2 (
         nx12903z23), .I3 (nx12903z25), .I4 (nx12903z24), .I5 (nx12903z19)) ;
         defparam ix12903z55292.INIT = 64'h9A4C2D3665B9D26C;
    (* HLUTNM = "LUT62_1_15" *)
    LUT4 ix42825z28456 (.O (nx42825z143), .I0 (\plaintext(20)  ), .I1 (nx37232z6
         ), .I2 (nx36230z5), .I3 (nx9305z5)) ;
         defparam ix42825z28456.INIT = 16'h6996;
    LUT6 ix12903z28451 (.O (nx12903z108), .I0 (\plaintext(36)  ), .I1 (
         \p_key_samp(45)  ), .I2 (nx37232z11), .I3 (px3635), .I4 (px3436), .I5 (
         px3197)) ;
         defparam ix12903z28451.INIT = 64'h6996966996696996;
    LUT6 ix12903z51430 (.O (px3197), .I0 (nx12903z40), .I1 (nx12903z42), .I2 (
         nx12903z43), .I3 (nx12903z44), .I4 (nx12903z45), .I5 (nx12903z47)) ;
         defparam ix12903z51430.INIT = 64'hA56A56A93C97C358;
    (* HLUTNM = "LUT62_1_13" *)
    LUT4 ix52909z39819 (.O (px3198), .I0 (\plaintext(36)  ), .I1 (nx37232z11), .I2 (
         px3635), .I3 (px3436)) ;
         defparam ix52909z39819.INIT = 16'h9669;
    LUT6 ix12903z28449 (.O (nx12903z106), .I0 (\plaintext(12)  ), .I1 (
         \p_key_samp(12)  ), .I2 (nx37232z4), .I3 (nx36230z3), .I4 (nx9305z3), .I5 (
         nx12903z107)) ;
         defparam ix12903z28449.INIT = 64'h6996966996696996;
    LUT6 ix12903z37853 (.O (nx12903z107), .I0 (nx12903z30), .I1 (nx12903z32), .I2 (
         nx12903z33), .I3 (nx12903z34), .I4 (nx12903z35), .I5 (nx12903z37)) ;
         defparam ix12903z37853.INIT = 64'h9672768B316D8E51;
    (* HLUTNM = "LUT62_1_14" *)
    LUT4 ix42825z39942 (.O (nx42825z156), .I0 (\plaintext(12)  ), .I1 (nx37232z4
         ), .I2 (nx36230z3), .I3 (nx9305z3)) ;
         defparam ix42825z39942.INIT = 16'h9669;
    (* HLUTNM = "LUT62_1_62" *)
    LUT4 ix54899z39819 (.O (px3202), .I0 (\plaintext(61)  ), .I1 (nx37232z2), .I2 (
         px3632), .I3 (px3392)) ;
         defparam ix54899z39819.INIT = 16'h9669;
    LUT6 ix12903z28436 (.O (nx12903z93), .I0 (\plaintext(11)  ), .I1 (
         \p_key_samp(11)  ), .I2 (nx16286z6), .I3 (nx13298z76), .I4 (nx12903z6)
         , .I5 (nx12903z94)) ;
         defparam ix12903z28436.INIT = 64'h6996966996696996;
    LUT6 ix12903z52527 (.O (nx12903z94), .I0 (nx12903z95), .I1 (nx12903z96), .I2 (
         nx12903z98), .I3 (nx12903z100), .I4 (nx12903z102), .I5 (nx12903z103)) ;
         defparam ix12903z52527.INIT = 64'h792C596A2A5DC7B0;
    LUT6 ix12903z39921 (.O (nx12903z103), .I0 (plaintext[2]), .I1 (
         \p_key_samp(61)  ), .I2 (nx40221z2), .I3 (px3674), .I4 (px3483), .I5 (
         px3206)) ;
         defparam ix12903z39921.INIT = 64'h9669699669969669;
    LUT6 ix32966z39748 (.O (px3206), .I0 (nx32966z3), .I1 (nx32966z4), .I2 (
         nx32966z5), .I3 (nx32966z6), .I4 (nx32966z8), .I5 (nx32966z10)) ;
         defparam ix32966z39748.INIT = 64'h96A6C3657A6D9621;
    (* HLUTNM = "LUT62_1_1" *)
    LUT4 ix54904z39819 (.O (px3207), .I0 (plaintext[2]), .I1 (nx40221z2), .I2 (
         px3674), .I3 (px3483)) ;
         defparam ix54904z39819.INIT = 16'h9669;
    LUT6 ix12903z28445 (.O (nx12903z102), .I0 (\plaintext(30)  ), .I1 (
         \p_key_samp(5)  ), .I2 (nx63157z44), .I3 (px3752), .I4 (px3523), .I5 (
         px3283)) ;
         defparam ix12903z28445.INIT = 64'h6996966996696996;
    LUT6 ix12903z28443 (.O (nx12903z100), .I0 (\plaintext(54)  ), .I1 (
         \p_key_samp(29)  ), .I2 (nx34235z34), .I3 (nx13298z15), .I4 (nx3326z5)
         , .I5 (nx12903z101)) ;
         defparam ix12903z28443.INIT = 64'h6996966996696996;
    LUT6 ix12903z36031 (.O (nx12903z101), .I0 (nx35956z7), .I1 (nx35956z5), .I2 (
         nx35956z3), .I3 (nx35956z10), .I4 (nx35956z9), .I5 (nx35956z8)) ;
         defparam ix12903z36031.INIT = 64'h8E3539C669CA8739;
    (* HLUTNM = "LUT62_1_10" *)
    LUT4 ix42825z39854 (.O (nx42825z41), .I0 (\plaintext(54)  ), .I1 (nx34235z34
         ), .I2 (nx13298z15), .I3 (nx3326z5)) ;
         defparam ix42825z39854.INIT = 16'h9669;
    LUT6 ix12903z39916 (.O (nx12903z98), .I0 (\plaintext(46)  ), .I1 (
         \p_key_samp(7)  ), .I2 (nx34235z37), .I3 (nx13298z13), .I4 (nx3326z8), 
         .I5 (nx12903z99)) ;
         defparam ix12903z39916.INIT = 64'h9669699669969669;
    LUT6 ix12903z27670 (.O (nx12903z99), .I0 (nx12903z52), .I1 (nx12903z53), .I2 (
         nx12903z54), .I3 (nx12903z56), .I4 (nx12903z57), .I5 (nx12903z59)) ;
         defparam ix12903z27670.INIT = 64'h69B869E599656692;
    (* HLUTNM = "LUT62_1_11" *)
    LUT4 ix42825z39828 (.O (nx42825z12), .I0 (\plaintext(46)  ), .I1 (nx34235z37
         ), .I2 (nx13298z13), .I3 (nx3326z8)) ;
         defparam ix42825z39828.INIT = 16'h9669;
    LUT6 ix12903z39914 (.O (nx12903z96), .I0 (\plaintext(62)  ), .I1 (
         \p_key_samp(55)  ), .I2 (nx37232z13), .I3 (nx36230z11), .I4 (nx9305z10)
         , .I5 (px3216)) ;
         defparam ix12903z39914.INIT = 64'h9669699669969669;
    LUT6 ix12903z41540 (.O (px3216), .I0 (nx12903z5), .I1 (nx12903z7), .I2 (
         nx12903z9), .I3 (nx12903z10), .I4 (nx12903z11), .I5 (nx12903z12)) ;
         defparam ix12903z41540.INIT = 64'h258B5B65563E9CC2;
    (* HLUTNM = "LUT62_1_12" *)
    LUT4 ix55901z39819 (.O (px3217), .I0 (\plaintext(62)  ), .I1 (nx37232z13), .I2 (
         nx36230z11), .I3 (nx9305z10)) ;
         defparam ix55901z39819.INIT = 16'h9669;
    LUT6 ix12903z28438 (.O (nx12903z95), .I0 (\plaintext(38)  ), .I1 (
         \p_key_samp(46)  ), .I2 (nx63157z36), .I3 (px3726), .I4 (px3582), .I5 (
         px3296)) ;
         defparam ix12903z28438.INIT = 64'h6996966996696996;
    (* HLUTNM = "LUT62_1_43" *)
    LUT4 ix42825z39825 (.O (nx42825z9), .I0 (\plaintext(11)  ), .I1 (nx16286z6)
         , .I2 (nx13298z76), .I3 (nx12903z6)) ;
         defparam ix42825z39825.INIT = 16'h9669;
    LUT6 ix12903z39900 (.O (nx12903z82), .I0 (plaintext[3]), .I1 (
         \p_key_samp(18)  ), .I2 (nx38222z2), .I3 (px3649), .I4 (px3405), .I5 (
         px3221)) ;
         defparam ix12903z39900.INIT = 64'h9669699669969669;
    LUT6 ix12903z27154 (.O (px3221), .I0 (nx12903z84), .I1 (nx12903z86), .I2 (
         nx12903z87), .I3 (nx12903z89), .I4 (nx12903z91), .I5 (nx12903z92)) ;
         defparam ix12903z27154.INIT = 64'h533EE9C0B9D0649E;
    (* HLUTNM = "LUT62_1_63" *)
    LUT4 ix56893z28344 (.O (px3222), .I0 (plaintext[3]), .I1 (nx38222z2), .I2 (
         px3649), .I3 (px3405)) ;
         defparam ix56893z28344.INIT = 16'h6996;
    LUT6 ix12903z28403 (.O (nx12903z60), .I0 (\plaintext(19)  ), .I1 (
         \p_key_samp(59)  ), .I2 (nx16286z9), .I3 (nx13298z72), .I4 (nx12903z8)
         , .I5 (nx12903z61)) ;
         defparam ix12903z28403.INIT = 64'h6996966996696996;
    LUT6 ix12903z51384 (.O (nx12903z61), .I0 (nx12903z62), .I1 (nx12903z64), .I2 (
         nx12903z66), .I3 (nx12903z68), .I4 (nx12903z70), .I5 (nx12903z80)) ;
         defparam ix12903z51384.INIT = 64'h552AB3C62CB5C35A;
    LUT6 ix12903z28423 (.O (nx12903z80), .I0 (\plaintext(26)  ), .I1 (
         \p_key_samp(58)  ), .I2 (nx45210z2), .I3 (px3716), .I4 (px3454), .I5 (
         px3226)) ;
         defparam ix12903z28423.INIT = 64'h6996966996696996;
    LUT6 ix12903z48126 (.O (px3226), .I0 (nx12903z30), .I1 (nx12903z32), .I2 (
         nx12903z33), .I3 (nx12903z34), .I4 (nx12903z35), .I5 (nx12903z37)) ;
         defparam ix12903z48126.INIT = 64'hD16E4E698A71B68C;
    (* HLUTNM = "LUT62_1_19" *)
    LUT4 ix56898z28344 (.O (px3227), .I0 (\plaintext(26)  ), .I1 (nx45210z2), .I2 (
         px3716), .I3 (px3454)) ;
         defparam ix56898z28344.INIT = 16'h6996;
    LUT6 ix12903z39888 (.O (nx12903z70), .I0 (\plaintext(34)  ), .I1 (
         \p_key_samp(44)  ), .I2 (nx41222z2), .I3 (px3688), .I4 (px3448), .I5 (
         px3229)) ;
         defparam ix12903z39888.INIT = 64'h9669699669969669;
    LUT6 ix12903z51412 (.O (px3229), .I0 (nx12903z72), .I1 (nx12903z73), .I2 (
         nx12903z74), .I3 (nx12903z75), .I4 (nx12903z76), .I5 (nx12903z78)) ;
         defparam ix12903z51412.INIT = 64'h6D5926B66983C36C;
    (* HLUTNM = "LUT62_1_20" *)
    LUT4 ix57888z28344 (.O (px3230), .I0 (\plaintext(34)  ), .I1 (nx41222z2), .I2 (
         px3688), .I3 (px3448)) ;
         defparam ix57888z28344.INIT = 16'h6996;
    LUT6 ix12903z39886 (.O (nx12903z68), .I0 (\plaintext(58)  ), .I1 (
         \p_key_samp(19)  ), .I2 (nx34235z18), .I3 (px3705), .I4 (px3460), .I5 (
         px3232)) ;
         defparam ix12903z39886.INIT = 64'h9669699669969669;
    LUT6 ix12903z16173 (.O (px3232), .I0 (nx12903z52), .I1 (nx12903z53), .I2 (
         nx12903z57), .I3 (nx12903z59), .I4 (nx12903z54), .I5 (nx12903z56)) ;
         defparam ix12903z16173.INIT = 64'h39D65AA8C63839C7;
    (* HLUTNM = "LUT62_1_26" *)
    LUT4 ix57891z39819 (.O (px3233), .I0 (\plaintext(58)  ), .I1 (nx34235z18), .I2 (
         px3705), .I3 (px3460)) ;
         defparam ix57891z39819.INIT = 16'h9669;
    LUT6 ix12903z28409 (.O (nx12903z66), .I0 (plaintext[6]), .I1 (
         \p_key_samp(41)  ), .I2 (nx44209z2), .I3 (px3702), .I4 (px3451), .I5 (
         px3235)) ;
         defparam ix12903z28409.INIT = 64'h6996966996696996;
    LUT6 ix12903z37530 (.O (px3235), .I0 (nx12903z10), .I1 (nx12903z9), .I2 (
         nx12903z12), .I3 (nx12903z7), .I4 (nx12903z5), .I5 (nx12903z11)) ;
         defparam ix12903z37530.INIT = 64'h943D62CA4FF08D36;
    (* HLUTNM = "LUT62_1_24" *)
    LUT4 ix57894z39819 (.O (px3236), .I0 (plaintext[6]), .I1 (nx44209z2), .I2 (
         px3702), .I3 (px3451)) ;
         defparam ix57894z39819.INIT = 16'h9669;
    LUT6 ix12903z28407 (.O (nx12903z64), .I0 (\plaintext(42)  ), .I1 (
         \p_key_samp(2)  ), .I2 (nx34235z15), .I3 (nx7313z4), .I4 (nx7312z3), .I5 (
         nx12903z65)) ;
         defparam ix12903z28407.INIT = 64'h6996966996696996;
    LUT6 ix12903z28926 (.O (nx12903z65), .I0 (nx35956z9), .I1 (nx35956z7), .I2 (
         nx35956z8), .I3 (nx35956z3), .I4 (nx35956z5), .I5 (nx35956z10)) ;
         defparam ix12903z28926.INIT = 64'hA13ECCC3D2256B9C;
    (* HLUTNM = "LUT62_1_23" *)
    LUT4 ix42825z28416 (.O (nx42825z86), .I0 (\plaintext(42)  ), .I1 (nx34235z15
         ), .I2 (nx7313z4), .I3 (nx7312z3)) ;
         defparam ix42825z28416.INIT = 16'h6996;
    LUT6 ix12903z39880 (.O (nx12903z62), .I0 (\plaintext(50)  ), .I1 (
         \p_key_samp(17)  ), .I2 (nx34235z13), .I3 (nx7313z10), .I4 (nx7312z7), 
         .I5 (nx12903z63)) ;
         defparam ix12903z39880.INIT = 64'h9669699669969669;
    LUT6 ix12903z23594 (.O (nx12903z63), .I0 (nx32966z3), .I1 (nx32966z5), .I2 (
         nx32966z6), .I3 (nx32966z4), .I4 (nx32966z10), .I5 (nx32966z8)) ;
         defparam ix12903z23594.INIT = 64'h49179671A6AD56CA;
    (* HLUTNM = "LUT62_1_25" *)
    LUT4 ix42825z28405 (.O (nx42825z72), .I0 (\plaintext(50)  ), .I1 (nx34235z13
         ), .I2 (nx7313z10), .I3 (nx7312z7)) ;
         defparam ix42825z28405.INIT = 16'h6996;
    (* HLUTNM = "LUT62_1_37" *)
    LUT4 ix42825z28402 (.O (nx42825z68), .I0 (\plaintext(19)  ), .I1 (nx16286z9)
         , .I2 (nx13298z72), .I3 (nx12903z8)) ;
         defparam ix42825z28402.INIT = 16'h6996;
    LUT6 ix12903z39832 (.O (nx12903z14), .I0 (\plaintext(35)  ), .I1 (
         \p_key_samp(42)  ), .I2 (nx39226z2), .I3 (px3652), .I4 (px3408), .I5 (
         px3245)) ;
         defparam ix12903z39832.INIT = 64'h9669699669969669;
    LUT6 ix12903z43918 (.O (px3245), .I0 (nx12903z16), .I1 (nx12903z26), .I2 (
         nx12903z28), .I3 (nx12903z38), .I4 (nx12903z48), .I5 (nx12903z50)) ;
         defparam ix12903z43918.INIT = 64'hE21D39D44DA2A65E;
    LUT6 ix12903z39868 (.O (nx12903z50), .I0 (\plaintext(40)  ), .I1 (
         \p_key_samp(57)  ), .I2 (nx39226z7), .I3 (nx24265z12), .I4 (nx5318z9), 
         .I5 (nx12903z51)) ;
         defparam ix12903z39868.INIT = 64'h9669699669969669;
    LUT6 ix12903z20151 (.O (nx12903z51), .I0 (nx12903z52), .I1 (nx12903z53), .I2 (
         nx12903z54), .I3 (nx12903z56), .I4 (nx12903z57), .I5 (nx12903z59)) ;
         defparam ix12903z20151.INIT = 64'h09A2F7BCB48D4963;
    LUT5 ix12903z28402 (.O (nx12903z59), .I0 (\plaintext(29)  ), .I1 (
         \p_key_samp(14)  ), .I2 (nx23267z2), .I3 (px3511), .I4 (px3321)) ;
         defparam ix12903z28402.INIT = 32'h96696996;
    LUT5 ix12903z28400 (.O (nx12903z57), .I0 (\plaintext(13)  ), .I1 (
         \p_key_samp(61)  ), .I2 (nx15291z29), .I3 (nx13298z29), .I4 (nx12903z58
         )) ;
         defparam ix12903z28400.INIT = 32'h96696996;
    LUT6 ix12903z24564 (.O (nx12903z58), .I0 (nx13298z2), .I1 (nx13298z22), .I2 (
         nx13298z36), .I3 (nx13298z47), .I4 (nx13298z59), .I5 (nx13298z69)) ;
         defparam ix12903z24564.INIT = 64'h3943677886A75A99;
    (* HLUTNM = "LUT62_1_51" *)
    LUT3 ix42825z1442 (.O (nx42825z26), .I0 (\plaintext(13)  ), .I1 (nx15291z29)
         , .I2 (nx13298z29)) ;
         defparam ix42825z1442.INIT = 8'h69;
    LUT5 ix12903z39874 (.O (nx12903z56), .I0 (\p_plaintext(63)  ), .I1 (
         \p_key_samp(55)  ), .I2 (nx29253z2), .I3 (px3565), .I4 (px3359)) ;
         defparam ix12903z39874.INIT = 32'h69969669;
    LUT5 ix12903z28397 (.O (nx12903z54), .I0 (\plaintext(21)  ), .I1 (
         \p_key_samp(62)  ), .I2 (nx15291z32), .I3 (nx13298z25), .I4 (nx12903z55
         )) ;
         defparam ix12903z28397.INIT = 32'h96696996;
    LUT6 ix12903z30450 (.O (nx12903z55), .I0 (nx7312z8), .I1 (nx7312z18), .I2 (
         nx7312z4), .I3 (nx7312z2), .I4 (nx7312z20), .I5 (nx7312z6)) ;
         defparam ix12903z30450.INIT = 64'hDA95876C2768719A;
    (* HLUTNM = "LUT62_1_50" *)
    LUT3 ix42825z1476 (.O (nx42825z15), .I0 (\plaintext(21)  ), .I1 (nx15291z32)
         , .I2 (nx13298z25)) ;
         defparam ix42825z1476.INIT = 8'h96;
    LUT5 ix12903z28396 (.O (nx12903z53), .I0 (\p_plaintext(37)  ), .I1 (
         \p_key_samp(29)  ), .I2 (px3745), .I3 (px3514), .I4 (px3315)) ;
         defparam ix12903z28396.INIT = 32'h96696996;
    LUT5 ix12903z28395 (.O (nx12903z52), .I0 (p_nbus_plaintext[63]), .I1 (
         \p_key_samp(23)  ), .I2 (nx63157z2), .I3 (px3724), .I4 (px3504)) ;
         defparam ix12903z28395.INIT = 32'h96696996;
    (* HLUTNM = "LUT62_1_31" *)
    LUT4 ix42825z39965 (.O (nx42825z190), .I0 (\plaintext(40)  ), .I1 (nx39226z7
         ), .I2 (nx24265z12), .I3 (nx5318z9)) ;
         defparam ix42825z39965.INIT = 16'h9669;
    LUT6 ix12903z28391 (.O (nx12903z48), .I0 (\plaintext(56)  ), .I1 (
         \p_key_samp(50)  ), .I2 (nx63157z20), .I3 (nx27254z2), .I4 (px3536), .I5 (
         px3330)) ;
         defparam ix12903z28391.INIT = 64'h6996966996696996;
    LUT6 ix12903z28381 (.O (nx12903z38), .I0 (\plaintext(24)  ), .I1 (
         \p_key_samp(25)  ), .I2 (nx39226z17), .I3 (px3657), .I4 (px3410), .I5 (
         px3261)) ;
         defparam ix12903z28381.INIT = 64'h6996966996696996;
    LUT6 ix12903z28430 (.O (px3261), .I0 (nx12903z40), .I1 (nx12903z42), .I2 (
         nx12903z43), .I3 (nx12903z44), .I4 (nx12903z45), .I5 (nx12903z47)) ;
         defparam ix12903z28430.INIT = 64'h9C61933D996669C6;
    (* HLUTNM = "LUT62_1_28" *)
    LUT4 ix60881z28344 (.O (px3262), .I0 (\plaintext(24)  ), .I1 (nx39226z17), .I2 (
         px3657), .I3 (px3410)) ;
         defparam ix60881z28344.INIT = 16'h6996;
    LUT6 ix12903z28371 (.O (nx12903z28), .I0 (plaintext[0]), .I1 (
         \p_key_samp(11)  ), .I2 (nx63157z28), .I3 (px3739), .I4 (px3506), .I5 (
         px3313)) ;
         defparam ix12903z28371.INIT = 64'h6996966996696996;
    LUT6 ix12903z28369 (.O (nx12903z26), .I0 (\plaintext(48)  ), .I1 (
         \p_key_samp(43)  ), .I2 (nx39226z4), .I3 (nx24265z7), .I4 (nx5318z6), .I5 (
         nx12903z27)) ;
         defparam ix12903z28369.INIT = 64'h6996966996696996;
    LUT6 ix12903z59586 (.O (nx12903z27), .I0 (nx32966z3), .I1 (nx32966z4), .I2 (
         nx32966z5), .I3 (nx32966z6), .I4 (nx32966z8), .I5 (nx32966z10)) ;
         defparam ix12903z59586.INIT = 64'hE79A54291675E386;
    LUT5 ix32966z28353 (.O (nx32966z10), .I0 (\plaintext(57)  ), .I1 (
         \p_key_samp(12)  ), .I2 (nx34235z21), .I3 (px3596), .I4 (px3307)) ;
         defparam ix32966z28353.INIT = 32'h96696996;
    LUT5 ix32966z28351 (.O (nx32966z8), .I0 (\plaintext(15)  ), .I1 (
         \p_key_samp(53)  ), .I2 (nx15291z18), .I3 (nx13298z54), .I4 (nx32966z9)
         ) ;
         defparam ix32966z28351.INIT = 32'h96696996;
    LUT6 ix32966z63762 (.O (nx32966z9), .I0 (nx3326z2), .I1 (nx3326z3), .I2 (
         nx3326z4), .I3 (nx3326z6), .I4 (nx3326z7), .I5 (nx3326z9)) ;
         defparam ix32966z63762.INIT = 64'h56298C178697F3E8;
    (* HLUTNM = "LUT62_1_52" *)
    LUT3 ix12903z1655 (.O (nx12903z252), .I0 (\plaintext(15)  ), .I1 (nx15291z18
         ), .I2 (nx13298z54)) ;
         defparam ix12903z1655.INIT = 8'h69;
    LUT5 ix32966z39824 (.O (nx32966z6), .I0 (\plaintext(23)  ), .I1 (
         \p_key_samp(63)  ), .I2 (nx15291z24), .I3 (nx13298z50), .I4 (nx32966z7)
         ) ;
         defparam ix32966z39824.INIT = 32'h69969669;
    LUT6 ix32966z13312 (.O (nx32966z7), .I0 (nx4319z2), .I1 (nx4319z4), .I2 (
         nx4319z6), .I3 (nx4319z7), .I4 (nx4319z8), .I5 (nx4319z9)) ;
         defparam ix32966z13312.INIT = 64'h394DC327A1972ED8;
    (* HLUTNM = "LUT62_1_53" *)
    LUT3 ix42825z1528 (.O (nx42825z75), .I0 (\plaintext(23)  ), .I1 (nx15291z24)
         , .I2 (nx13298z50)) ;
         defparam ix42825z1528.INIT = 8'h96;
    LUT5 ix32966z28348 (.O (nx32966z5), .I0 (\p_plaintext(39)  ), .I1 (
         \p_key_samp(5)  ), .I2 (px3781), .I3 (px3559), .I4 (px3353)) ;
         defparam ix32966z28348.INIT = 32'h96696996;
    LUT5 ix32966z39822 (.O (nx32966z4), .I0 (\plaintext(31)  ), .I1 (
         \p_key_samp(38)  ), .I2 (nx28253z2), .I3 (px3562), .I4 (px3373)) ;
         defparam ix32966z39822.INIT = 32'h69969669;
    LUT5 ix32966z28346 (.O (nx32966z3), .I0 (\plaintext(7)  ), .I1 (
         \p_key_samp(7)  ), .I2 (nx34235z6), .I3 (px3587), .I4 (px3304)) ;
         defparam ix32966z28346.INIT = 32'h96696996;
    (* HLUTNM = "LUT62_1_30" *)
    LUT4 ix42825z28487 (.O (nx42825z186), .I0 (\plaintext(48)  ), .I1 (nx39226z4
         ), .I2 (nx24265z7), .I3 (nx5318z6)) ;
         defparam ix42825z28487.INIT = 16'h6996;
    LUT6 ix12903z28359 (.O (nx12903z16), .I0 (\plaintext(32)  ), .I1 (
         \p_key_samp(60)  ), .I2 (nx39226z15), .I3 (px3665), .I4 (px3421), .I5 (
         px3278)) ;
         defparam ix12903z28359.INIT = 64'h6996966996696996;
    LUT6 ix12903z48535 (.O (px3278), .I0 (nx12903z18), .I1 (nx12903z19), .I2 (
         nx12903z21), .I3 (nx12903z23), .I4 (nx12903z24), .I5 (nx12903z25)) ;
         defparam ix12903z48535.INIT = 64'hB1494BB45AB6B865;
    (* HLUTNM = "LUT62_1_27" *)
    LUT4 ix61885z28344 (.O (px3279), .I0 (\plaintext(32)  ), .I1 (nx39226z15), .I2 (
         px3665), .I3 (px3421)) ;
         defparam ix61885z28344.INIT = 16'h6996;
    (* HLUTNM = "LUT62_1_64" *)
    LUT4 ix62873z39819 (.O (px3280), .I0 (\plaintext(35)  ), .I1 (nx39226z2), .I2 (
         px3652), .I3 (px3408)) ;
         defparam ix62873z39819.INIT = 16'h9669;
    LUT6 ix12903z13859 (.O (px3281), .I0 (nx12903z91), .I1 (nx12903z87), .I2 (
         nx12903z92), .I3 (nx12903z86), .I4 (nx12903z84), .I5 (nx12903z89)) ;
         defparam ix12903z13859.INIT = 64'hBA5157AC473C306B;
    LUT6 ix12903z28432 (.O (nx12903z89), .I0 (\plaintext(30)  ), .I1 (
         \p_key_samp(54)  ), .I2 (nx63157z44), .I3 (px3752), .I4 (px3523), .I5 (
         px3283)) ;
         defparam ix12903z28432.INIT = 64'h6996966996696996;
    LUT6 ix12903z48128 (.O (px3283), .I0 (nx12903z18), .I1 (nx12903z21), .I2 (
         nx12903z23), .I3 (nx12903z25), .I4 (nx12903z24), .I5 (nx12903z19)) ;
         defparam ix12903z48128.INIT = 64'hB6878B788C78B685;
    LUT5 ix12903z39837 (.O (nx12903z19), .I0 (\plaintext(51)  ), .I1 (
         \p_key_samp(1)  ), .I2 (nx25263z8), .I3 (nx24265z37), .I4 (nx12903z20)
         ) ;
         defparam ix12903z39837.INIT = 32'h69969669;
    LUT6 ix12903z31469 (.O (nx12903z20), .I0 (nx11304z2), .I1 (nx11304z4), .I2 (
         nx11304z5), .I3 (nx11304z7), .I4 (nx11304z8), .I5 (nx11304z9)) ;
         defparam ix12903z31469.INIT = 64'h4B911E2D946E75B8;
    (* HLUTNM = "LUT62_1_48" *)
    LUT3 ix42825z1583 (.O (nx42825z151), .I0 (\plaintext(51)  ), .I1 (nx25263z8)
         , .I2 (nx24265z37)) ;
         defparam ix42825z1583.INIT = 8'h96;
    LUT5 ix12903z28367 (.O (nx12903z24), .I0 (\plaintext(27)  ), .I1 (
         \p_key_samp(42)  ), .I2 (nx36228z2), .I3 (px3615), .I4 (px3425)) ;
         defparam ix12903z28367.INIT = 32'h96696996;
    LUT5 ix12903z39843 (.O (nx12903z25), .I0 (\plaintext(59)  ), .I1 (
         \p_key_samp(3)  ), .I2 (nx27254z4), .I3 (px3546), .I4 (px3338)) ;
         defparam ix12903z39843.INIT = 32'h69969669;
    LUT5 ix12903z28366 (.O (nx12903z23), .I0 (plaintext[5]), .I1 (
         \p_key_samp(25)  ), .I2 (nx27254z7), .I3 (px3543), .I4 (px3341)) ;
         defparam ix12903z28366.INIT = 32'h96696996;
    LUT5 ix12903z28364 (.O (nx12903z21), .I0 (\plaintext(43)  ), .I1 (
         \p_key_samp(49)  ), .I2 (nx25263z6), .I3 (nx24265z26), .I4 (nx12903z22)
         ) ;
         defparam ix12903z28364.INIT = 32'h96696996;
    LUT6 ix12903z37528 (.O (nx12903z22), .I0 (nx337z9), .I1 (nx337z3), .I2 (
         nx337z8), .I3 (nx337z2), .I4 (nx337z5), .I5 (nx337z7)) ;
         defparam ix12903z37528.INIT = 64'hEC21C33E789E8D61;
    (* HLUTNM = "LUT62_1_41" *)
    LUT3 ix42825z1579 (.O (nx42825z146), .I0 (\plaintext(43)  ), .I1 (nx25263z6)
         , .I2 (nx24265z26)) ;
         defparam ix42825z1579.INIT = 8'h96;
    LUT5 ix12903z39836 (.O (nx12903z18), .I0 (\plaintext(35)  ), .I1 (
         \p_key_samp(59)  ), .I2 (nx39226z2), .I3 (px3652), .I4 (px3408)) ;
         defparam ix12903z39836.INIT = 32'h69969669;
    (* HLUTNM = "LUT62_1_7" *)
    LUT4 ix63874z28344 (.O (px3294), .I0 (\plaintext(30)  ), .I1 (nx63157z44), .I2 (
         px3752), .I3 (px3523)) ;
         defparam ix63874z28344.INIT = 16'h6996;
    LUT6 ix12903z28427 (.O (nx12903z84), .I0 (\plaintext(38)  ), .I1 (
         \p_key_samp(21)  ), .I2 (nx63157z36), .I3 (px3726), .I4 (px3582), .I5 (
         px3296)) ;
         defparam ix12903z28427.INIT = 64'h6996966996696996;
    LUT6 ix12903z39240 (.O (px3296), .I0 (nx12903z72), .I1 (nx12903z73), .I2 (
         nx12903z74), .I3 (nx12903z75), .I4 (nx12903z76), .I5 (nx12903z78)) ;
         defparam ix12903z39240.INIT = 64'hA6C949357C6A93D2;
    LUT5 ix12903z28421 (.O (nx12903z78), .I0 (\plaintext(49)  ), .I1 (
         \p_key_samp(27)  ), .I2 (nx34235z4), .I3 (nx13298z62), .I4 (nx12903z79)
         ) ;
         defparam ix12903z28421.INIT = 32'h96696996;
    LUT6 ix12903z28482 (.O (nx12903z79), .I0 (nx11304z2), .I1 (nx11304z4), .I2 (
         nx11304z5), .I3 (nx11304z7), .I4 (nx11304z8), .I5 (nx11304z9)) ;
         defparam ix12903z28482.INIT = 64'hD10CB46BAA7969D2;
    (* HLUTNM = "LUT62_1_42" *)
    LUT3 ix42825z1567 (.O (nx42825z128), .I0 (\plaintext(49)  ), .I1 (nx34235z4)
         , .I2 (nx13298z62)) ;
         defparam ix42825z1567.INIT = 8'h96;
    LUT5 ix12903z39894 (.O (nx12903z76), .I0 (\plaintext(41)  ), .I1 (
         \p_key_samp(41)  ), .I2 (nx34235z8), .I3 (nx13298z65), .I4 (nx12903z77)
         ) ;
         defparam ix12903z39894.INIT = 32'h69969669;
    LUT6 ix12903z55060 (.O (nx12903z77), .I0 (nx9305z2), .I1 (nx9305z4), .I2 (
         nx9305z6), .I3 (nx9305z7), .I4 (nx9305z8), .I5 (nx9305z9)) ;
         defparam ix12903z55060.INIT = 64'h57896596E453D1A6;
    (* HLUTNM = "LUT62_1_49" *)
    LUT3 ix42825z1525 (.O (nx42825z132), .I0 (\plaintext(41)  ), .I1 (nx34235z8)
         , .I2 (nx13298z65)) ;
         defparam ix42825z1525.INIT = 8'h69;
    LUT5 ix12903z28418 (.O (nx12903z75), .I0 (\plaintext(7)  ), .I1 (
         \p_key_samp(58)  ), .I2 (nx34235z6), .I3 (px3587), .I4 (px3304)) ;
         defparam ix12903z28418.INIT = 32'h96696996;
    LUT6 ix334z40647 (.O (px3304), .I0 (nx13298z2), .I1 (nx13298z22), .I2 (
         nx13298z36), .I3 (nx13298z47), .I4 (nx13298z59), .I5 (nx13298z69)) ;
         defparam ix334z40647.INIT = 64'h43C67898A77999A5;
    (* HLUTNM = "LUT62_1_33" *)
    LUT3 ix335z1464 (.O (px3305), .I0 (\plaintext(7)  ), .I1 (nx34235z6), .I2 (
         px3587)) ;
         defparam ix335z1464.INIT = 8'h96;
    LUT5 ix12903z28417 (.O (nx12903z74), .I0 (\plaintext(57)  ), .I1 (
         \p_key_samp(34)  ), .I2 (nx34235z21), .I3 (px3596), .I4 (px3307)) ;
         defparam ix12903z28417.INIT = 32'h96696996;
    LUT6 ix337z59898 (.O (px3307), .I0 (nx337z2), .I1 (nx337z3), .I2 (nx337z5), 
         .I3 (nx337z7), .I4 (nx337z8), .I5 (nx337z9)) ;
         defparam ix337z59898.INIT = 64'hE15E99691E91E4D8;
    (* HLUTNM = "LUT62_1_34" *)
    LUT3 ix338z1464 (.O (px3308), .I0 (\plaintext(57)  ), .I1 (nx34235z21), .I2 (
         px3596)) ;
         defparam ix338z1464.INIT = 8'h96;
    LUT5 ix12903z28416 (.O (nx12903z73), .I0 (\plaintext(25)  ), .I1 (
         \p_key_samp(9)  ), .I2 (nx34235z31), .I3 (px3590), .I4 (px3335)) ;
         defparam ix12903z28416.INIT = 32'h96696996;
    LUT5 ix12903z28415 (.O (nx12903z72), .I0 (\plaintext(33)  ), .I1 (
         \p_key_samp(44)  ), .I2 (nx34235z10), .I3 (px3584), .I4 (px3332)) ;
         defparam ix12903z28415.INIT = 32'h96696996;
    (* HLUTNM = "LUT62_1_8" *)
    LUT4 ix1328z28344 (.O (px3311), .I0 (\plaintext(38)  ), .I1 (nx63157z36), .I2 (
         px3726), .I3 (px3582)) ;
         defparam ix1328z28344.INIT = 16'h6996;
    LUT6 ix12903z28429 (.O (nx12903z86), .I0 (plaintext[0]), .I1 (
         \p_key_samp(23)  ), .I2 (nx63157z28), .I3 (px3739), .I4 (px3506), .I5 (
         px3313)) ;
         defparam ix12903z28429.INIT = 64'h6996966996696996;
    LUT6 ix12903z60504 (.O (px3313), .I0 (nx12903z30), .I1 (nx12903z32), .I2 (
         nx12903z33), .I3 (nx12903z34), .I4 (nx12903z35), .I5 (nx12903z37)) ;
         defparam ix12903z60504.INIT = 64'h662868B71CD9E71A;
    LUT5 ix12903z28380 (.O (nx12903z37), .I0 (\p_plaintext(37)  ), .I1 (
         \p_key_samp(21)  ), .I2 (px3745), .I3 (px3514), .I4 (px3315)) ;
         defparam ix12903z28380.INIT = 32'h96696996;
    LUT6 ix1332z27325 (.O (px3315), .I0 (nx3326z2), .I1 (nx3326z3), .I2 (
         nx3326z4), .I3 (nx3326z6), .I4 (nx3326z7), .I5 (nx3326z9)) ;
         defparam ix1332z27325.INIT = 64'h3C69D23C8B64659B;
    (* HLUTNM = "LUT62_1_35" *)
    LUT3 ix1333z1419 (.O (px3316), .I0 (\p_plaintext(37)  ), .I1 (px3745), .I2 (
         px3514)) ;
         defparam ix1333z1419.INIT = 8'h69;
    LUT5 ix12903z39853 (.O (nx12903z35), .I0 (\plaintext(45)  ), .I1 (
         \p_key_samp(22)  ), .I2 (nx16289z7), .I3 (nx7312z12), .I4 (nx12903z36)
         ) ;
         defparam ix12903z39853.INIT = 32'h69969669;
    LUT6 ix12903z15248 (.O (nx12903z36), .I0 (nx4319z4), .I1 (nx4319z7), .I2 (
         nx4319z6), .I3 (nx4319z2), .I4 (nx4319z8), .I5 (nx4319z9)) ;
         defparam ix12903z15248.INIT = 64'h964EE1994BB4364B;
    (* HLUTNM = "LUT62_1_47" *)
    LUT3 ix42825z1557 (.O (nx42825z113), .I0 (\plaintext(45)  ), .I1 (nx16289z7)
         , .I2 (nx7312z12)) ;
         defparam ix42825z1557.INIT = 8'h96;
    LUT5 ix12903z28377 (.O (nx12903z34), .I0 (\plaintext(29)  ), .I1 (
         \p_key_samp(28)  ), .I2 (nx23267z2), .I3 (px3511), .I4 (px3321)) ;
         defparam ix12903z28377.INIT = 32'h96696996;
    LUT6 ix2325z20403 (.O (px3321), .I0 (nx337z2), .I1 (nx337z3), .I2 (nx337z5)
         , .I3 (nx337z7), .I4 (nx337z8), .I5 (nx337z9)) ;
         defparam ix2325z20403.INIT = 64'h7227B55EACD84A91;
    (* HLUTNM = "LUT62_1_36" *)
    LUT3 ix2326z1464 (.O (px3322), .I0 (\plaintext(29)  ), .I1 (nx23267z2), .I2 (
         px3511)) ;
         defparam ix2326z1464.INIT = 8'h96;
    LUT5 ix12903z28376 (.O (nx12903z33), .I0 (plaintext[3]), .I1 (
         \p_key_samp(46)  ), .I2 (nx38222z2), .I3 (px3649), .I4 (px3405)) ;
         defparam ix12903z28376.INIT = 32'h96696996;
    LUT5 ix12903z39850 (.O (nx12903z32), .I0 (\plaintext(61)  ), .I1 (
         \p_key_samp(4)  ), .I2 (nx37232z2), .I3 (px3632), .I4 (px3392)) ;
         defparam ix12903z39850.INIT = 32'h69969669;
    LUT5 ix12903z39848 (.O (nx12903z30), .I0 (\plaintext(53)  ), .I1 (
         \p_key_samp(31)  ), .I2 (nx16289z10), .I3 (nx7312z17), .I4 (nx12903z31)
         ) ;
         defparam ix12903z39848.INIT = 32'h69969669;
    LUT6 ix12903z39947 (.O (nx12903z31), .I0 (nx5318z2), .I1 (nx5318z3), .I2 (
         nx5318z5), .I3 (nx5318z8), .I4 (nx5318z4), .I5 (nx5318z7)) ;
         defparam ix12903z39947.INIT = 64'hAAD525A5562996CB;
    (* HLUTNM = "LUT62_1_46" *)
    LUT3 ix42825z1509 (.O (nx42825z110), .I0 (\plaintext(53)  ), .I1 (nx16289z10
         ), .I2 (nx7312z17)) ;
         defparam ix42825z1509.INIT = 8'h69;
    (* HLUTNM = "LUT62_1_6" *)
    LUT4 ix2332z28344 (.O (px3328), .I0 (plaintext[0]), .I1 (nx63157z28), .I2 (
         px3739), .I3 (px3506)) ;
         defparam ix2332z28344.INIT = 16'h6996;
    LUT6 ix12903z28435 (.O (nx12903z92), .I0 (\plaintext(56)  ), .I1 (
         \p_key_samp(28)  ), .I2 (nx63157z20), .I3 (nx27254z2), .I4 (px3536), .I5 (
         px3330)) ;
         defparam ix12903z28435.INIT = 64'h6996966996696996;
    LUT6 ix12903z12684 (.O (px3330), .I0 (nx35956z3), .I1 (nx35956z5), .I2 (
         nx35956z7), .I3 (nx35956z8), .I4 (nx35956z9), .I5 (nx35956z10)) ;
         defparam ix12903z12684.INIT = 64'hA63C59A35B962C3A;
    LUT5 ix35956z28353 (.O (nx35956z10), .I0 (\plaintext(33)  ), .I1 (
         \p_key_samp(2)  ), .I2 (nx34235z10), .I3 (px3584), .I4 (px3332)) ;
         defparam ix35956z28353.INIT = 32'h96696996;
    LUT6 ix3323z29144 (.O (px3332), .I0 (nx7312z6), .I1 (nx7312z20), .I2 (
         nx7312z2), .I3 (nx7312z8), .I4 (nx7312z4), .I5 (nx7312z18)) ;
         defparam ix3323z29144.INIT = 64'h4BB8B1C3B4496CB6;
    (* HLUTNM = "LUT62_1_59" *)
    LUT3 ix3324z1464 (.O (px3333), .I0 (\plaintext(33)  ), .I1 (nx34235z10), .I2 (
         px3584)) ;
         defparam ix3324z1464.INIT = 8'h96;
    LUT5 ix35956z28352 (.O (nx35956z9), .I0 (\plaintext(25)  ), .I1 (
         \p_key_samp(11)  ), .I2 (nx34235z31), .I3 (px3590), .I4 (px3335)) ;
         defparam ix35956z28352.INIT = 32'h96696996;
    LUT6 ix3326z39864 (.O (px3335), .I0 (nx3326z2), .I1 (nx3326z3), .I2 (
         nx3326z4), .I3 (nx3326z6), .I4 (nx3326z7), .I5 (nx3326z9)) ;
         defparam ix3326z39864.INIT = 64'h956796896A969696;
    (* HLUTNM = "LUT62_1_58" *)
    LUT3 ix42825z1518 (.O (nx42825z60), .I0 (\plaintext(25)  ), .I1 (nx34235z31)
         , .I2 (px3590)) ;
         defparam ix42825z1518.INIT = 8'h96;
    LUT5 ix35956z39826 (.O (nx35956z8), .I0 (\plaintext(59)  ), .I1 (
         \p_key_samp(60)  ), .I2 (nx27254z4), .I3 (px3546), .I4 (px3338)) ;
         defparam ix35956z39826.INIT = 32'h69969669;
    LUT6 ix3329z51039 (.O (px3338), .I0 (nx9305z6), .I1 (nx9305z2), .I2 (
         nx9305z8), .I3 (nx9305z4), .I4 (nx9305z9), .I5 (nx9305z7)) ;
         defparam ix3329z51039.INIT = 64'hD2662DD26D8AC23D;
    (* HLUTNM = "LUT62_1_60" *)
    LUT3 ix42825z1463 (.O (nx42825z50), .I0 (\plaintext(59)  ), .I1 (nx27254z4)
         , .I2 (px3546)) ;
         defparam ix42825z1463.INIT = 8'h69;
    LUT5 ix35956z28350 (.O (nx35956z7), .I0 (plaintext[5]), .I1 (
         \p_key_samp(33)  ), .I2 (nx27254z7), .I3 (px3543), .I4 (px3341)) ;
         defparam ix35956z28350.INIT = 32'h96696996;
    LUT6 ix4319z43150 (.O (px3341), .I0 (nx4319z2), .I1 (nx4319z4), .I2 (
         nx4319z6), .I3 (nx4319z7), .I4 (nx4319z8), .I5 (nx4319z9)) ;
         defparam ix4319z43150.INIT = 64'h5A35963915CEA36C;
    (* HLUTNM = "LUT62_1_57" *)
    LUT3 ix4320z1419 (.O (px3342), .I0 (plaintext[5]), .I1 (nx27254z7), .I2 (
         px3543)) ;
         defparam ix4320z1419.INIT = 8'h69;
    LUT5 ix35956z39823 (.O (nx35956z5), .I0 (\plaintext(17)  ), .I1 (
         \p_key_samp(26)  ), .I2 (nx27254z11), .I3 (nx13298z9), .I4 (nx35956z6)
         ) ;
         defparam ix35956z39823.INIT = 32'h69969669;
    LUT6 ix35956z39373 (.O (nx35956z6), .I0 (nx5318z2), .I1 (nx5318z3), .I2 (
         nx5318z5), .I3 (nx5318z8), .I4 (nx5318z4), .I5 (nx5318z7)) ;
         defparam ix35956z39373.INIT = 64'h369C96C36B9594A6;
    (* HLUTNM = "LUT62_1_45" *)
    LUT3 ix42825z1512 (.O (nx42825z54), .I0 (\plaintext(17)  ), .I1 (nx27254z11)
         , .I2 (nx13298z9)) ;
         defparam ix42825z1512.INIT = 8'h96;
    LUT5 ix35956z28346 (.O (nx35956z3), .I0 (\plaintext(9)  ), .I1 (
         \p_key_samp(51)  ), .I2 (nx27254z9), .I3 (nx13298z5), .I4 (nx35956z4)
         ) ;
         defparam ix35956z28346.INIT = 32'h96696996;
    LUT6 ix35956z15185 (.O (nx35956z4), .I0 (nx13298z2), .I1 (nx13298z22), .I2 (
         nx13298z36), .I3 (nx13298z47), .I4 (nx13298z59), .I5 (nx13298z69)) ;
         defparam ix35956z15185.INIT = 64'h5A99E95E91E1362C;
    (* HLUTNM = "LUT62_1_40" *)
    LUT3 ix42825z1505 (.O (nx42825z47), .I0 (\plaintext(9)  ), .I1 (nx27254z9), 
         .I2 (nx13298z5)) ;
         defparam ix42825z1505.INIT = 8'h96;
    (* HLUTNM = "LUT62_1_5" *)
    LUT4 ix4327z28344 (.O (px3349), .I0 (\plaintext(56)  ), .I1 (nx63157z20), .I2 (
         nx27254z2), .I3 (px3536)) ;
         defparam ix4327z28344.INIT = 16'h6996;
    LUT6 ix12903z39905 (.O (nx12903z87), .I0 (\plaintext(14)  ), .I1 (
         \p_key_samp(4)  ), .I2 (nx63157z12), .I3 (nx37234z7), .I4 (nx11304z6), 
         .I5 (nx12903z88)) ;
         defparam ix12903z39905.INIT = 64'h9669699669969669;
    LUT6 ix12903z27697 (.O (nx12903z88), .I0 (nx12903z40), .I1 (nx12903z42), .I2 (
         nx12903z43), .I3 (nx12903z44), .I4 (nx12903z45), .I5 (nx12903z47)) ;
         defparam ix12903z27697.INIT = 64'h2EF8CB96510766B8;
    LUT5 ix12903z28390 (.O (nx12903z47), .I0 (\p_plaintext(39)  ), .I1 (
         \p_key_samp(30)  ), .I2 (px3781), .I3 (px3559), .I4 (px3353)) ;
         defparam ix12903z28390.INIT = 32'h96696996;
    LUT6 ix5318z36612 (.O (px3353), .I0 (nx5318z2), .I1 (nx5318z3), .I2 (
         nx5318z4), .I3 (nx5318z5), .I4 (nx5318z7), .I5 (nx5318z8)) ;
         defparam ix5318z36612.INIT = 64'h49B0355EB65E89E2;
    (* HLUTNM = "LUT62_1_54" *)
    LUT3 ix5319z1464 (.O (px3354), .I0 (\p_plaintext(39)  ), .I1 (px3781), .I2 (
         px3559)) ;
         defparam ix5319z1464.INIT = 8'h96;
    LUT5 ix12903z28388 (.O (nx12903z45), .I0 (\plaintext(47)  ), .I1 (
         \p_key_samp(20)  ), .I2 (nx15291z12), .I3 (nx13298z46), .I4 (nx12903z46
         )) ;
         defparam ix12903z28388.INIT = 32'h96696996;
    LUT6 ix12903z8196 (.O (nx12903z46), .I0 (nx9305z2), .I1 (nx9305z4), .I2 (
         nx9305z6), .I3 (nx9305z7), .I4 (nx9305z8), .I5 (nx9305z9)) ;
         defparam ix12903z8196.INIT = 64'h3CA5C35A36691AB5;
    (* HLUTNM = "LUT62_1_39" *)
    LUT3 ix12903z2249 (.O (nx12903z453), .I0 (\plaintext(47)  ), .I1 (nx15291z12
         ), .I2 (nx13298z46)) ;
         defparam ix12903z2249.INIT = 8'h96;
    LUT5 ix12903z39862 (.O (nx12903z44), .I0 (\p_plaintext(63)  ), .I1 (
         \p_key_samp(39)  ), .I2 (nx29253z2), .I3 (px3565), .I4 (px3359)) ;
         defparam ix12903z39862.INIT = 32'h69969669;
    LUT6 ix5324z40936 (.O (px3359), .I0 (nx4319z2), .I1 (nx4319z4), .I2 (
         nx4319z6), .I3 (nx4319z7), .I4 (nx4319z8), .I5 (nx4319z9)) ;
         defparam ix5324z40936.INIT = 64'h74A9A17AD31C9AC6;
    LUT5 ix4319z39827 (.O (nx4319z9), .I0 (\plaintext(60)  ), .I1 (
         \p_key_samp(51)  ), .I2 (nx36228z10), .I3 (px3623), .I4 (px3439)) ;
         defparam ix4319z39827.INIT = 32'h69969669;
    LUT5 ix4319z28351 (.O (nx4319z8), .I0 (\plaintext(34)  ), .I1 (
         \p_key_samp(2)  ), .I2 (nx41222z2), .I3 (px3688), .I4 (px3448)) ;
         defparam ix4319z28351.INIT = 32'h96696996;
    LUT5 ix4319z28350 (.O (nx4319z7), .I0 (plaintext[4]), .I1 (\p_key_samp(41)  
         ), .I2 (nx36228z6), .I3 (px3626), .I4 (px3433)) ;
         defparam ix4319z28350.INIT = 32'h96696996;
    LUT5 ix4319z28349 (.O (nx4319z6), .I0 (\plaintext(26)  ), .I1 (
         \p_key_samp(1)  ), .I2 (nx45210z2), .I3 (px3716), .I4 (px3454)) ;
         defparam ix4319z28349.INIT = 32'h96696996;
    LUT5 ix4319z39822 (.O (nx4319z4), .I0 (\plaintext(18)  ), .I1 (
         \p_key_samp(19)  ), .I2 (nx29253z8), .I3 (nx24265z20), .I4 (nx4319z5)
         ) ;
         defparam ix4319z39822.INIT = 32'h69969669;
    LUT6 ix4319z14738 (.O (nx4319z5), .I0 (nx24265z13), .I1 (nx24265z15), .I2 (
         nx24265z25), .I3 (nx24265z35), .I4 (nx24265z36), .I5 (nx24265z2)) ;
         defparam ix4319z14738.INIT = 64'h55CAEA93A539346C;
    (* HLUTNM = "LUT62_1_77" *)
    LUT3 ix12903z1828 (.O (nx12903z472), .I0 (\plaintext(18)  ), .I1 (nx29253z8)
         , .I2 (nx24265z20)) ;
         defparam ix12903z1828.INIT = 8'h69;
    LUT5 ix4319z39820 (.O (nx4319z2), .I0 (\plaintext(10)  ), .I1 (
         \p_key_samp(34)  ), .I2 (nx29253z10), .I3 (nx24265z23), .I4 (nx4319z3)
         ) ;
         defparam ix4319z39820.INIT = 32'h69969669;
    LUT6 ix4319z41670 (.O (nx4319z3), .I0 (nx13298z41), .I1 (nx13298z42), .I2 (
         nx13298z40), .I3 (nx13298z38), .I4 (nx13298z45), .I5 (nx13298z44)) ;
         defparam ix4319z41670.INIT = 64'h3B1CC3E458679DA2;
    (* HLUTNM = "LUT62_1_79" *)
    LUT3 ix12903z1832 (.O (nx12903z477), .I0 (\plaintext(10)  ), .I1 (nx29253z10
         ), .I2 (nx24265z23)) ;
         defparam ix12903z1832.INIT = 8'h69;
    (* HLUTNM = "LUT62_1_56" *)
    LUT3 ix12903z1824 (.O (nx12903z467), .I0 (\p_plaintext(63)  ), .I1 (
         nx29253z2), .I2 (px3565)) ;
         defparam ix12903z1824.INIT = 8'h69;
    LUT5 ix12903z28386 (.O (nx12903z43), .I0 (p_nbus_plaintext[63]), .I1 (
         \p_key_samp(45)  ), .I2 (nx63157z2), .I3 (px3724), .I4 (px3504)) ;
         defparam ix12903z28386.INIT = 32'h96696996;
    LUT5 ix12903z39860 (.O (nx12903z42), .I0 (\plaintext(31)  ), .I1 (
         \p_key_samp(54)  ), .I2 (nx28253z2), .I3 (px3562), .I4 (px3373)) ;
         defparam ix12903z39860.INIT = 32'h69969669;
    LUT6 ix7312z46716 (.O (px3373), .I0 (nx7312z2), .I1 (nx7312z4), .I2 (
         nx7312z6), .I3 (nx7312z8), .I4 (nx7312z18), .I5 (nx7312z20)) ;
         defparam ix7312z46716.INIT = 64'hBCCB4B741661B15A;
    (* HLUTNM = "LUT62_1_55" *)
    LUT3 ix7313z1464 (.O (px3374), .I0 (\plaintext(31)  ), .I1 (nx28253z2), .I2 (
         px3562)) ;
         defparam ix7313z1464.INIT = 8'h96;
    LUT5 ix12903z39858 (.O (nx12903z40), .I0 (\plaintext(55)  ), .I1 (
         \p_key_samp(13)  ), .I2 (nx15291z8), .I3 (nx13298z39), .I4 (nx12903z41)
         ) ;
         defparam ix12903z39858.INIT = 32'h69969669;
    LUT6 ix12903z13072 (.O (nx12903z41), .I0 (nx337z2), .I1 (nx337z3), .I2 (
         nx337z5), .I3 (nx337z7), .I4 (nx337z8), .I5 (nx337z9)) ;
         defparam ix12903z13072.INIT = 64'h2BC5963AC6392DC6;
    LUT5 ix337z28352 (.O (nx337z9), .I0 (\plaintext(24)  ), .I1 (
         \p_key_samp(58)  ), .I2 (nx39226z17), .I3 (px3657), .I4 (px3410)) ;
         defparam ix337z28352.INIT = 32'h96696996;
    LUT5 ix337z39826 (.O (nx337z8), .I0 (\plaintext(58)  ), .I1 (
         \p_key_samp(44)  ), .I2 (nx34235z18), .I3 (px3705), .I4 (px3460)) ;
         defparam ix337z39826.INIT = 32'h69969669;
    LUT5 ix337z28350 (.O (nx337z7), .I0 (\plaintext(32)  ), .I1 (
         \p_key_samp(49)  ), .I2 (nx39226z15), .I3 (px3665), .I4 (px3421)) ;
         defparam ix337z28350.INIT = 32'h96696996;
    LUT5 ix337z28348 (.O (nx337z5), .I0 (\plaintext(8)  ), .I1 (\p_key_samp(35)  
         ), .I2 (nx34235z25), .I3 (nx24265z31), .I4 (nx337z6)) ;
         defparam ix337z28348.INIT = 32'h96696996;
    LUT6 ix337z20818 (.O (nx337z6), .I0 (nx7312z10), .I1 (nx7312z11), .I2 (
         nx7312z13), .I3 (nx7312z14), .I4 (nx7312z15), .I5 (nx7312z16)) ;
         defparam ix337z20818.INIT = 64'h4B9C9E74B0D64C2B;
    (* HLUTNM = "LUT62_1_38" *)
    LUT3 ix12903z1833 (.O (nx12903z425), .I0 (\plaintext(8)  ), .I1 (nx34235z25)
         , .I2 (nx24265z31)) ;
         defparam ix12903z1833.INIT = 8'h96;
    LUT5 ix337z39821 (.O (nx337z3), .I0 (\plaintext(16)  ), .I1 (
         \p_key_samp(10)  ), .I2 (nx34235z28), .I3 (nx24265z33), .I4 (nx337z4)
         ) ;
         defparam ix337z39821.INIT = 32'h69969669;
    LUT6 ix337z28654 (.O (nx337z4), .I0 (nx13298z61), .I1 (nx13298z63), .I2 (
         nx13298z64), .I3 (nx13298z66), .I4 (nx13298z67), .I5 (nx13298z68)) ;
         defparam ix337z28654.INIT = 64'h8BA9743C95566AC9;
    (* HLUTNM = "LUT62_1_78" *)
    LUT3 ix12903z1830 (.O (nx12903z421), .I0 (\plaintext(16)  ), .I1 (nx34235z28
         ), .I2 (nx24265z33)) ;
         defparam ix12903z1830.INIT = 8'h96;
    LUT5 ix337z39820 (.O (nx337z2), .I0 (plaintext[6]), .I1 (\p_key_samp(17)  )
         , .I2 (nx44209z2), .I3 (px3702), .I4 (px3451)) ;
         defparam ix337z39820.INIT = 32'h69969669;
    (* HLUTNM = "LUT62_1_44" *)
    LUT3 ix12903z1827 (.O (nx12903z417), .I0 (\plaintext(55)  ), .I1 (nx15291z8)
         , .I2 (nx13298z39)) ;
         defparam ix12903z1827.INIT = 8'h96;
    (* HLUTNM = "LUT62_1_9" *)
    LUT4 ix12903z40163 (.O (nx12903z392), .I0 (\plaintext(14)  ), .I1 (
         nx63157z12), .I2 (nx37234z7), .I3 (nx11304z6)) ;
         defparam ix12903z40163.INIT = 16'h9669;
    LUT6 ix12903z28434 (.O (nx12903z91), .I0 (\plaintext(22)  ), .I1 (
         \p_key_samp(14)  ), .I2 (nx63157z4), .I3 (nx37234z3), .I4 (nx11304z3), 
         .I5 (nx12903z4)) ;
         defparam ix12903z28434.INIT = 64'h6996966996696996;
    LUT6 ix12903z46702 (.O (nx12903z4), .I0 (nx12903z5), .I1 (nx12903z7), .I2 (
         nx12903z9), .I3 (nx12903z10), .I4 (nx12903z11), .I5 (nx12903z12)) ;
         defparam ix12903z46702.INIT = 64'hC39C4E172EDAB149;
    LUT5 ix12903z39830 (.O (nx12903z12), .I0 (\plaintext(61)  ), .I1 (
         \p_key_samp(36)  ), .I2 (nx37232z2), .I3 (px3632), .I4 (px3392)) ;
         defparam ix12903z39830.INIT = 32'h69969669;
    LUT6 ix9305z23469 (.O (px3392), .I0 (nx9305z2), .I1 (nx9305z4), .I2 (
         nx9305z6), .I3 (nx9305z7), .I4 (nx9305z8), .I5 (nx9305z9)) ;
         defparam ix9305z23469.INIT = 64'h7A43297CA53C568B;
    LUT5 ix9305z39827 (.O (nx9305z9), .I0 (\plaintext(62)  ), .I1 (
         \p_key_samp(39)  ), .I2 (nx37232z13), .I3 (nx36230z11), .I4 (nx9305z10)
         ) ;
         defparam ix9305z39827.INIT = 32'h69969669;
    LUT5 ix9305z39826 (.O (nx9305z8), .I0 (\plaintext(36)  ), .I1 (
         \p_key_samp(13)  ), .I2 (nx37232z11), .I3 (px3635), .I4 (px3436)) ;
         defparam ix9305z39826.INIT = 32'h69969669;
    LUT5 ix9305z39825 (.O (nx9305z7), .I0 (\plaintext(28)  ), .I1 (
         \p_key_samp(63)  ), .I2 (nx37232z9), .I3 (px3638), .I4 (px3442)) ;
         defparam ix9305z39825.INIT = 32'h69969669;
    LUT5 ix9305z39824 (.O (nx9305z6), .I0 (plaintext[2]), .I1 (\p_key_samp(7)  )
         , .I2 (nx40221z2), .I3 (px3674), .I4 (px3483)) ;
         defparam ix9305z39824.INIT = 32'h69969669;
    LUT5 ix9305z28347 (.O (nx9305z4), .I0 (\plaintext(20)  ), .I1 (
         \p_key_samp(46)  ), .I2 (nx37232z6), .I3 (nx36230z5), .I4 (nx9305z5)) ;
         defparam ix9305z28347.INIT = 32'h96696996;
    LUT6 ix9305z47756 (.O (nx9305z5), .I0 (nx24265z2), .I1 (nx24265z13), .I2 (
         nx24265z15), .I3 (nx24265z25), .I4 (nx24265z35), .I5 (nx24265z36)) ;
         defparam ix9305z47756.INIT = 64'hB60D489B68D3B566;
    (* HLUTNM = "LUT62_1_80" *)
    LUT3 ix12903z1860 (.O (nx12903z457), .I0 (\plaintext(20)  ), .I1 (nx37232z6)
         , .I2 (nx36230z5)) ;
         defparam ix12903z1860.INIT = 8'h96;
    LUT5 ix9305z39820 (.O (nx9305z2), .I0 (\plaintext(12)  ), .I1 (
         \p_key_samp(45)  ), .I2 (nx37232z4), .I3 (nx36230z3), .I4 (nx9305z3)) ;
         defparam ix9305z39820.INIT = 32'h69969669;
    LUT6 ix9305z20192 (.O (nx9305z3), .I0 (nx7312z10), .I1 (nx7312z11), .I2 (
         nx7312z14), .I3 (nx7312z13), .I4 (nx7312z15), .I5 (nx7312z16)) ;
         defparam ix9305z20192.INIT = 64'h94B2A34D1BC749BC;
    (* HLUTNM = "LUT62_1_76" *)
    LUT3 ix12903z1818 (.O (nx12903z460), .I0 (\plaintext(12)  ), .I1 (nx37232z4)
         , .I2 (nx36230z3)) ;
         defparam ix12903z1818.INIT = 8'h69;
    (* HLUTNM = "LUT62_1_62" *)
    LUT3 ix11302z1419 (.O (px3403), .I0 (\plaintext(61)  ), .I1 (nx37232z2), .I2 (
         px3632)) ;
         defparam ix11302z1419.INIT = 8'h69;
    LUT5 ix12903z28354 (.O (nx12903z11), .I0 (plaintext[3]), .I1 (
         \p_key_samp(57)  ), .I2 (nx38222z2), .I3 (px3649), .I4 (px3405)) ;
         defparam ix12903z28354.INIT = 32'h96696996;
    LUT6 ix11304z8859 (.O (px3405), .I0 (nx11304z2), .I1 (nx11304z4), .I2 (
         nx11304z5), .I3 (nx11304z7), .I4 (nx11304z8), .I5 (nx11304z9)) ;
         defparam ix11304z8859.INIT = 64'hAD5A668B83451D79;
    (* HLUTNM = "LUT62_1_63" *)
    LUT3 ix11305z1464 (.O (px3406), .I0 (plaintext[3]), .I1 (nx38222z2), .I2 (
         px3649)) ;
         defparam ix11305z1464.INIT = 8'h96;
    LUT5 ix12903z39828 (.O (nx12903z10), .I0 (\plaintext(35)  ), .I1 (
         \p_key_samp(18)  ), .I2 (nx39226z2), .I3 (px3652), .I4 (px3408)) ;
         defparam ix12903z39828.INIT = 32'h69969669;
    LUT6 ix11307z45433 (.O (px3408), .I0 (nx5318z2), .I1 (nx5318z3), .I2 (
         nx5318z5), .I3 (nx5318z8), .I4 (nx5318z4), .I5 (nx5318z7)) ;
         defparam ix11307z45433.INIT = 64'h2D5653E8B298AC57;
    LUT5 ix5318z28350 (.O (nx5318z7), .I0 (\plaintext(24)  ), .I1 (
         \p_key_samp(60)  ), .I2 (nx39226z17), .I3 (px3657), .I4 (px3410)) ;
         defparam ix5318z28350.INIT = 32'h96696996;
    LUT6 ix12296z18616 (.O (px3410), .I0 (nx13298z38), .I1 (nx13298z40), .I2 (
         nx13298z41), .I3 (nx13298z42), .I4 (nx13298z44), .I5 (nx13298z45)) ;
         defparam ix12296z18616.INIT = 64'h96967C961EE14396;
    (* HLUTNM = "LUT62_1_66" *)
    LUT3 ix12297z1464 (.O (px3411), .I0 (\plaintext(24)  ), .I1 (nx39226z17), .I2 (
         px3657)) ;
         defparam ix12297z1464.INIT = 8'h96;
    LUT5 ix5318z28347 (.O (nx5318z4), .I0 (\plaintext(56)  ), .I1 (
         \p_key_samp(18)  ), .I2 (nx63157z20), .I3 (nx27254z2), .I4 (px3536)) ;
         defparam ix5318z28347.INIT = 32'h96696996;
    LUT5 ix5318z39826 (.O (nx5318z8), .I0 (\plaintext(40)  ), .I1 (
         \p_key_samp(25)  ), .I2 (nx39226z7), .I3 (nx24265z12), .I4 (nx5318z9)
         ) ;
         defparam ix5318z39826.INIT = 32'h69969669;
    LUT6 ix5318z27205 (.O (nx5318z9), .I0 (nx13298z24), .I1 (nx13298z26), .I2 (
         nx13298z28), .I3 (nx13298z30), .I4 (nx13298z32), .I5 (nx13298z34)) ;
         defparam ix5318z27205.INIT = 64'hE19E5A072CCB651B;
    (* HLUTNM = "LUT62_1_74" *)
    LUT3 ix12903z1760 (.O (nx12903z388), .I0 (\plaintext(40)  ), .I1 (nx39226z7)
         , .I2 (nx24265z12)) ;
         defparam ix12903z1760.INIT = 8'h69;
    LUT5 ix5318z28348 (.O (nx5318z5), .I0 (\plaintext(48)  ), .I1 (
         \p_key_samp(11)  ), .I2 (nx39226z4), .I3 (nx24265z7), .I4 (nx5318z6)) ;
         defparam ix5318z28348.INIT = 32'h96696996;
    LUT6 ix5318z29186 (.O (nx5318z6), .I0 (nx13298z57), .I1 (nx13298z55), .I2 (
         nx13298z58), .I3 (nx13298z49), .I4 (nx13298z53), .I5 (nx13298z51)) ;
         defparam ix5318z29186.INIT = 64'h49DAB32986316CDB;
    (* HLUTNM = "LUT62_1_75" *)
    LUT3 ix12903z1802 (.O (nx12903z381), .I0 (\plaintext(48)  ), .I1 (nx39226z4)
         , .I2 (nx24265z7)) ;
         defparam ix12903z1802.INIT = 8'h96;
    LUT5 ix5318z28346 (.O (nx5318z3), .I0 (plaintext[0]), .I1 (\p_key_samp(42)  
         ), .I2 (nx63157z28), .I3 (px3739), .I4 (px3506)) ;
         defparam ix5318z28346.INIT = 32'h96696996;
    LUT5 ix5318z28345 (.O (nx5318z2), .I0 (\plaintext(32)  ), .I1 (
         \p_key_samp(59)  ), .I2 (nx39226z15), .I3 (px3665), .I4 (px3421)) ;
         defparam ix5318z28345.INIT = 32'h96696996;
    LUT6 ix13294z43901 (.O (px3421), .I0 (nx24265z2), .I1 (nx24265z36), .I2 (
         nx24265z15), .I3 (nx24265z25), .I4 (nx24265z35), .I5 (nx24265z13)) ;
         defparam ix13294z43901.INIT = 64'hB44B19B485B6A65B;
    (* HLUTNM = "LUT62_1_81" *)
    LUT3 ix13295z1464 (.O (px3422), .I0 (\plaintext(32)  ), .I1 (nx39226z15), .I2 (
         px3665)) ;
         defparam ix13295z1464.INIT = 8'h96;
    (* HLUTNM = "LUT62_1_64" *)
    LUT3 ix12903z2088 (.O (nx12903z377), .I0 (\plaintext(35)  ), .I1 (nx39226z2)
         , .I2 (px3652)) ;
         defparam ix12903z2088.INIT = 8'h69;
    LUT5 ix12903z28352 (.O (nx12903z9), .I0 (\plaintext(27)  ), .I1 (
         \p_key_samp(17)  ), .I2 (nx36228z2), .I3 (px3615), .I4 (px3425)) ;
         defparam ix12903z28352.INIT = 32'h96696996;
    LUT6 ix13298z12779 (.O (px3425), .I0 (nx13298z2), .I1 (nx13298z22), .I2 (
         nx13298z36), .I3 (nx13298z47), .I4 (nx13298z59), .I5 (nx13298z69)) ;
         defparam ix13298z12779.INIT = 64'h99A55E16E16E2CC9;
    LUT5 ix13298z39888 (.O (nx13298z69), .I0 (\plaintext(44)  ), .I1 (
         \p_key_samp(6)  ), .I2 (nx36228z4), .I3 (nx15291z38), .I4 (nx13298z70)
         ) ;
         defparam ix13298z39888.INIT = 32'h69969669;
    LUT6 ix13298z39823 (.O (nx13298z70), .I0 (nx13298z71), .I1 (nx13298z73), .I2 (
         nx13298z74), .I3 (nx13298z75), .I4 (nx13298z77), .I5 (nx13298z78)) ;
         defparam ix13298z39823.INIT = 64'hC62D2DD278999627;
    (* HLUTNM = "LUT62_1_92" *)
    LUT3 ix42825z1490 (.O (nx42825z31), .I0 (\plaintext(44)  ), .I1 (nx36228z4)
         , .I2 (nx15291z38)) ;
         defparam ix42825z1490.INIT = 8'h96;
    LUT5 ix13298z39878 (.O (nx13298z59), .I0 (\plaintext(52)  ), .I1 (
         \p_key_samp(15)  ), .I2 (nx36228z8), .I3 (nx15291z36), .I4 (nx13298z60)
         ) ;
         defparam ix13298z39878.INIT = 32'h69969669;
    LUT6 ix13298z19640 (.O (nx13298z60), .I0 (nx13298z61), .I1 (nx13298z63), .I2 (
         nx13298z64), .I3 (nx13298z66), .I4 (nx13298z67), .I5 (nx13298z68)) ;
         defparam ix13298z19640.INIT = 64'hAC1BB86547B4475A;
    (* HLUTNM = "LUT62_1_93" *)
    LUT3 ix42825z1496 (.O (nx42825z37), .I0 (\plaintext(52)  ), .I1 (nx36228z8)
         , .I2 (nx15291z36)) ;
         defparam ix42825z1496.INIT = 8'h96;
    LUT5 ix13298z28391 (.O (nx13298z47), .I0 (plaintext[4]), .I1 (
         \p_key_samp(30)  ), .I2 (nx36228z6), .I3 (px3626), .I4 (px3433)) ;
         defparam ix13298z28391.INIT = 32'h96696996;
    LUT6 ix13298z28418 (.O (px3433), .I0 (nx13298z49), .I1 (nx13298z51), .I2 (
         nx13298z53), .I3 (nx13298z55), .I4 (nx13298z57), .I5 (nx13298z58)) ;
         defparam ix13298z28418.INIT = 64'h66787989D1AE69B0;
    (* HLUTNM = "LUT62_1_82" *)
    LUT3 ix14294z1464 (.O (px3434), .I0 (plaintext[4]), .I1 (nx36228z6), .I2 (
         px3626)) ;
         defparam ix14294z1464.INIT = 8'h96;
    LUT5 ix13298z39855 (.O (nx13298z36), .I0 (\plaintext(36)  ), .I1 (
         \p_key_samp(5)  ), .I2 (nx37232z11), .I3 (px3635), .I4 (px3436)) ;
         defparam ix13298z39855.INIT = 32'h69969669;
    LUT6 ix13298z39803 (.O (px3436), .I0 (nx13298z38), .I1 (nx13298z40), .I2 (
         nx13298z41), .I3 (nx13298z42), .I4 (nx13298z44), .I5 (nx13298z45)) ;
         defparam ix13298z39803.INIT = 64'h59B466CB668B9634;
    (* HLUTNM = "LUT62_1_83" *)
    LUT3 ix14297z1419 (.O (px3437), .I0 (\plaintext(36)  ), .I1 (nx37232z11), .I2 (
         px3635)) ;
         defparam ix14297z1419.INIT = 8'h69;
    LUT5 ix13298z39841 (.O (nx13298z22), .I0 (\plaintext(60)  ), .I1 (
         \p_key_samp(53)  ), .I2 (nx36228z10), .I3 (px3623), .I4 (px3439)) ;
         defparam ix13298z39841.INIT = 32'h69969669;
    LUT6 ix13298z40565 (.O (px3439), .I0 (nx13298z24), .I1 (nx13298z26), .I2 (
         nx13298z28), .I3 (nx13298z30), .I4 (nx13298z32), .I5 (nx13298z34)) ;
         defparam ix13298z40565.INIT = 64'h931CE66946D3993C;
    (* HLUTNM = "LUT62_1_84" *)
    LUT3 ix15287z1419 (.O (px3440), .I0 (\plaintext(60)  ), .I1 (nx36228z10), .I2 (
         px3623)) ;
         defparam ix15287z1419.INIT = 8'h69;
    LUT5 ix13298z39820 (.O (nx13298z2), .I0 (\plaintext(28)  ), .I1 (
         \p_key_samp(12)  ), .I2 (nx37232z9), .I3 (px3638), .I4 (px3442)) ;
         defparam ix13298z39820.INIT = 32'h69969669;
    LUT6 ix13298z60719 (.O (px3442), .I0 (nx13298z4), .I1 (nx13298z6), .I2 (
         nx13298z7), .I3 (nx13298z8), .I4 (nx13298z10), .I5 (nx13298z20)) ;
         defparam ix13298z60719.INIT = 64'h29EBD69017D6E80B;
    (* HLUTNM = "LUT62_1_85" *)
    LUT3 ix15290z1419 (.O (px3443), .I0 (\plaintext(28)  ), .I1 (nx37232z9), .I2 (
         px3638)) ;
         defparam ix15290z1419.INIT = 8'h69;
    (* HLUTNM = "LUT62_1_61" *)
    LUT3 ix15291z1419 (.O (px3444), .I0 (\plaintext(27)  ), .I1 (nx36228z2), .I2 (
         px3615)) ;
         defparam ix15291z1419.INIT = 8'h69;
    LUT5 ix12903z28350 (.O (nx12903z7), .I0 (\plaintext(19)  ), .I1 (
         \p_key_samp(35)  ), .I2 (nx16286z9), .I3 (nx13298z72), .I4 (nx12903z8)
         ) ;
         defparam ix12903z28350.INIT = 32'h96696996;
    LUT6 ix12903z16752 (.O (nx12903z8), .I0 (nx7312z2), .I1 (nx7312z4), .I2 (
         nx7312z6), .I3 (nx7312z8), .I4 (nx7312z18), .I5 (nx7312z20)) ;
         defparam ix12903z16752.INIT = 64'hD947A9B82CB23C47;
    LUT5 ix7312z28363 (.O (nx7312z20), .I0 (\plaintext(34)  ), .I1 (
         \p_key_samp(43)  ), .I2 (nx41222z2), .I3 (px3688), .I4 (px3448)) ;
         defparam ix7312z28363.INIT = 32'h96696996;
    LUT6 ix7312z58980 (.O (px3448), .I0 (nx13298z61), .I1 (nx13298z63), .I2 (
         nx13298z64), .I3 (nx13298z66), .I4 (nx13298z67), .I5 (nx13298z68)) ;
         defparam ix7312z58980.INIT = 64'h3DC296788937E12E;
    (* HLUTNM = "LUT62_1_73" *)
    LUT3 ix12903z1759 (.O (nx12903z331), .I0 (\plaintext(34)  ), .I1 (nx41222z2)
         , .I2 (px3688)) ;
         defparam ix12903z1759.INIT = 8'h96;
    LUT5 ix7312z39836 (.O (nx7312z18), .I0 (plaintext[6]), .I1 (\p_key_samp(9)  
         ), .I2 (nx44209z2), .I3 (px3702), .I4 (px3451)) ;
         defparam ix7312z39836.INIT = 32'h69969669;
    LUT6 ix7312z41367 (.O (px3451), .I0 (nx13298z71), .I1 (nx13298z75), .I2 (
         nx13298z77), .I3 (nx13298z73), .I4 (nx13298z78), .I5 (nx13298z74)) ;
         defparam ix7312z41367.INIT = 64'h6A3D559CA25C9C63;
    (* HLUTNM = "LUT62_1_86" *)
    LUT3 ix16286z1419 (.O (px3452), .I0 (plaintext[6]), .I1 (nx44209z2), .I2 (
         px3702)) ;
         defparam ix16286z1419.INIT = 8'h69;
    LUT5 ix7312z28351 (.O (nx7312z8), .I0 (\plaintext(26)  ), .I1 (
         \p_key_samp(26)  ), .I2 (nx45210z2), .I3 (px3716), .I4 (px3454)) ;
         defparam ix7312z28351.INIT = 32'h96696996;
    LUT6 ix7312z56940 (.O (px3454), .I0 (nx7312z10), .I1 (nx7312z11), .I2 (
         nx7312z13), .I3 (nx7312z14), .I4 (nx7312z15), .I5 (nx7312z16)) ;
         defparam ix7312z56940.INIT = 64'hD23938ED25BCD942;
    (* HLUTNM = "LUT62_1_87" *)
    LUT3 ix16289z1464 (.O (px3455), .I0 (\plaintext(26)  ), .I1 (nx45210z2), .I2 (
         px3716)) ;
         defparam ix16289z1464.INIT = 8'h96;
    LUT5 ix7312z28349 (.O (nx7312z6), .I0 (\plaintext(50)  ), .I1 (
         \p_key_samp(52)  ), .I2 (nx34235z13), .I3 (nx7313z10), .I4 (nx7312z7)
         ) ;
         defparam ix7312z28349.INIT = 32'h96696996;
    LUT6 ix7312z26078 (.O (nx7312z7), .I0 (nx13298z57), .I1 (nx13298z58), .I2 (
         nx13298z49), .I3 (nx13298z55), .I4 (nx13298z53), .I5 (nx13298z51)) ;
         defparam ix7312z26078.INIT = 64'hB84D166B9FE060B6;
    (* HLUTNM = "LUT62_1_70" *)
    LUT3 ix12903z1748 (.O (nx12903z373), .I0 (\plaintext(50)  ), .I1 (nx34235z13
         ), .I2 (nx7313z10)) ;
         defparam ix12903z1748.INIT = 8'h69;
    LUT5 ix7312z39822 (.O (nx7312z4), .I0 (\plaintext(58)  ), .I1 (
         \p_key_samp(50)  ), .I2 (nx34235z18), .I3 (px3705), .I4 (px3460)) ;
         defparam ix7312z39822.INIT = 32'h69969669;
    LUT6 ix7312z15040 (.O (px3460), .I0 (nx13298z32), .I1 (nx13298z34), .I2 (
         nx13298z24), .I3 (nx13298z28), .I4 (nx13298z26), .I5 (nx13298z30)) ;
         defparam ix7312z15040.INIT = 64'h3C87DA68C369359A;
    (* HLUTNM = "LUT62_1_72" *)
    LUT3 ix12903z1755 (.O (nx12903z327), .I0 (\plaintext(58)  ), .I1 (nx34235z18
         ), .I2 (px3705)) ;
         defparam ix12903z1755.INIT = 8'h96;
    LUT5 ix7312z28345 (.O (nx7312z2), .I0 (\plaintext(42)  ), .I1 (
         \p_key_samp(33)  ), .I2 (nx34235z15), .I3 (nx7313z4), .I4 (nx7312z3)) ;
         defparam ix7312z28345.INIT = 32'h96696996;
    LUT6 ix7312z55113 (.O (nx7312z3), .I0 (nx13298z10), .I1 (nx13298z7), .I2 (
         nx13298z6), .I3 (nx13298z4), .I4 (nx13298z8), .I5 (nx13298z20)) ;
         defparam ix7312z55113.INIT = 64'hCCC3A13E6B9CD225;
    (* HLUTNM = "LUT62_1_71" *)
    LUT3 ix12903z1752 (.O (nx12903z322), .I0 (\plaintext(42)  ), .I1 (nx34235z15
         ), .I2 (nx7313z4)) ;
         defparam ix12903z1752.INIT = 8'h96;
    (* HLUTNM = "LUT62_1_37" *)
    LUT3 ix12903z1749 (.O (nx12903z319), .I0 (\plaintext(19)  ), .I1 (nx16286z9)
         , .I2 (nx13298z72)) ;
         defparam ix12903z1749.INIT = 8'h96;
    LUT5 ix12903z39823 (.O (nx12903z5), .I0 (\plaintext(11)  ), .I1 (
         \p_key_samp(50)  ), .I2 (nx16286z6), .I3 (nx13298z76), .I4 (nx12903z6)
         ) ;
         defparam ix12903z39823.INIT = 32'h69969669;
    LUT6 ix12903z13561 (.O (nx12903z6), .I0 (nx3326z2), .I1 (nx3326z3), .I2 (
         nx3326z4), .I3 (nx3326z6), .I4 (nx3326z7), .I5 (nx3326z9)) ;
         defparam ix12903z13561.INIT = 64'hB31DC4A61C5A2FD2;
    LUT5 ix3326z28352 (.O (nx3326z9), .I0 (\plaintext(38)  ), .I1 (
         \p_key_samp(14)  ), .I2 (nx63157z36), .I3 (px3726), .I4 (px3582)) ;
         defparam ix3326z28352.INIT = 32'h96696996;
    LUT5 ix3326z39825 (.O (nx3326z7), .I0 (\plaintext(46)  ), .I1 (
         \p_key_samp(4)  ), .I2 (nx34235z37), .I3 (nx13298z13), .I4 (nx3326z8)
         ) ;
         defparam ix3326z39825.INIT = 32'h69969669;
    LUT6 ix3326z35987 (.O (nx3326z8), .I0 (nx13298z24), .I1 (nx13298z26), .I2 (
         nx13298z28), .I3 (nx13298z30), .I4 (nx13298z32), .I5 (nx13298z34)) ;
         defparam ix3326z35987.INIT = 64'hC7263CD17855876A;
    LUT4 ix13298z39853 (.O (nx13298z34), .I0 (\p_plaintext(37)  ), .I1 (
         \p_key_samp(62)  ), .I2 (px3745), .I3 (px3514)) ;
         defparam ix13298z39853.INIT = 16'h9669;
    LUT4 ix13298z39851 (.O (nx13298z32), .I0 (p_nbus_plaintext[63]), .I1 (
         \p_key_samp(20)  ), .I2 (nx63157z2), .I3 (px3724)) ;
         defparam ix13298z39851.INIT = 16'h9669;
    LUT4 ix13298z28374 (.O (nx13298z30), .I0 (\plaintext(29)  ), .I1 (
         \p_key_samp(47)  ), .I2 (nx23267z2), .I3 (px3511)) ;
         defparam ix13298z28374.INIT = 16'h6996;
    LUT4 ix13298z39847 (.O (nx13298z28), .I0 (\plaintext(13)  ), .I1 (
         \p_key_samp(29)  ), .I2 (nx15291z29), .I3 (nx13298z29)) ;
         defparam ix13298z39847.INIT = 16'h9669;
    LUT6 ix13298z47064 (.O (nx13298z29), .I0 (nx15291z3), .I1 (nx15291z13), .I2 (
         nx15291z15), .I3 (nx15291z25), .I4 (nx15291z35), .I5 (nx15291z37)) ;
         defparam ix13298z47064.INIT = 64'h5B6CAD42C636B299;
    (* HLUTNM = "LUT62_1_81" *)
    LUT2 ix12903z1605 (.O (nx12903z310), .I0 (\plaintext(13)  ), .I1 (nx15291z29
         )) ;
         defparam ix12903z1605.INIT = 4'h9;
    LUT4 ix13298z39845 (.O (nx13298z26), .I0 (\p_plaintext(63)  ), .I1 (
         \p_key_samp(23)  ), .I2 (nx29253z2), .I3 (px3565)) ;
         defparam ix13298z39845.INIT = 16'h9669;
    LUT4 ix13298z28368 (.O (nx13298z24), .I0 (\plaintext(21)  ), .I1 (
         \p_key_samp(30)  ), .I2 (nx15291z32), .I3 (nx13298z25)) ;
         defparam ix13298z28368.INIT = 16'h6996;
    LUT6 ix13298z28046 (.O (nx13298z25), .I0 (nx7313z3), .I1 (nx7313z5), .I2 (
         nx7313z6), .I3 (nx7313z8), .I4 (nx7313z9), .I5 (nx7313z11)) ;
         defparam ix13298z28046.INIT = 64'hE952266D979C6853;
    (* HLUTNM = "LUT62_1_80" *)
    LUT2 ix12903z1599 (.O (nx12903z307), .I0 (\plaintext(21)  ), .I1 (nx15291z32
         )) ;
         defparam ix12903z1599.INIT = 4'h6;
    (* HLUTNM = "LUT62_1_68" *)
    LUT3 ix12903z1695 (.O (nx12903z304), .I0 (\plaintext(46)  ), .I1 (nx34235z37
         ), .I2 (nx13298z13)) ;
         defparam ix12903z1695.INIT = 8'h69;
    LUT5 ix3326z39824 (.O (nx3326z6), .I0 (plaintext[2]), .I1 (\p_key_samp(29)  
         ), .I2 (nx40221z2), .I3 (px3674), .I4 (px3483)) ;
         defparam ix3326z39824.INIT = 32'h69969669;
    LUT6 ix19278z4493 (.O (px3483), .I0 (nx13298z49), .I1 (nx13298z51), .I2 (
         nx13298z53), .I3 (nx13298z55), .I4 (nx13298z57), .I5 (nx13298z58)) ;
         defparam ix19278z4493.INIT = 64'hAE45533C57B80C6B;
    LUT4 ix13298z28402 (.O (nx13298z58), .I0 (\p_plaintext(39)  ), .I1 (
         \p_key_samp(38)  ), .I2 (px3781), .I3 (px3559)) ;
         defparam ix13298z28402.INIT = 16'h6996;
    LUT4 ix13298z28401 (.O (nx13298z57), .I0 (\plaintext(31)  ), .I1 (
         \p_key_samp(6)  ), .I2 (nx28253z2), .I3 (px3562)) ;
         defparam ix13298z28401.INIT = 16'h6996;
    LUT4 ix13298z28399 (.O (nx13298z55), .I0 (\plaintext(7)  ), .I1 (
         \p_key_samp(4)  ), .I2 (nx34235z6), .I3 (px3587)) ;
         defparam ix13298z28399.INIT = 16'h6996;
    LUT4 ix13298z39872 (.O (nx13298z53), .I0 (\plaintext(15)  ), .I1 (
         \p_key_samp(21)  ), .I2 (nx15291z18), .I3 (nx13298z54)) ;
         defparam ix13298z39872.INIT = 16'h9669;
    LUT6 ix13298z24576 (.O (nx13298z54), .I0 (nx13298z14), .I1 (nx13298z18), .I2 (
         nx13298z17), .I3 (nx13298z12), .I4 (nx13298z19), .I5 (nx13298z16)) ;
         defparam ix13298z24576.INIT = 64'h96CD3D53C5325AA8;
    LUT4 ix13298z28395 (.O (nx13298z51), .I0 (\plaintext(57)  ), .I1 (
         \p_key_samp(45)  ), .I2 (nx34235z21), .I3 (px3596)) ;
         defparam ix13298z28395.INIT = 16'h6996;
    LUT4 ix13298z28393 (.O (nx13298z49), .I0 (\plaintext(23)  ), .I1 (
         \p_key_samp(31)  ), .I2 (nx15291z24), .I3 (nx13298z50)) ;
         defparam ix13298z28393.INIT = 16'h6996;
    LUT6 ix13298z3789 (.O (nx13298z50), .I0 (nx24265z17), .I1 (nx24265z19), .I2 (
         nx24265z18), .I3 (nx24265z22), .I4 (nx24265z21), .I5 (nx24265z24)) ;
         defparam ix13298z3789.INIT = 64'h5F96B4C293A60979;
    (* HLUTNM = "LUT62_1_72" *)
    LUT2 ix12903z1532 (.O (nx12903z223), .I0 (\plaintext(23)  ), .I1 (nx15291z24
         )) ;
         defparam ix12903z1532.INIT = 4'h9;
    (* HLUTNM = "LUT62_1_67" *)
    LUT3 ix12903z1624 (.O (nx12903z218), .I0 (plaintext[2]), .I1 (nx40221z2), .I2 (
         px3674)) ;
         defparam ix12903z1624.INIT = 8'h69;
    LUT5 ix3326z39822 (.O (nx3326z4), .I0 (\plaintext(54)  ), .I1 (
         \p_key_samp(62)  ), .I2 (nx34235z34), .I3 (nx13298z15), .I4 (nx3326z5)
         ) ;
         defparam ix3326z39822.INIT = 32'h69969669;
    LUT6 ix3326z13048 (.O (nx3326z5), .I0 (nx13298z7), .I1 (nx13298z4), .I2 (
         nx13298z8), .I3 (nx13298z6), .I4 (nx13298z20), .I5 (nx13298z10)) ;
         defparam ix3326z13048.INIT = 64'h2B96D12ED2392DD2;
    (* HLUTNM = "LUT62_1_69" *)
    LUT3 ix12903z1706 (.O (nx12903z261), .I0 (\plaintext(54)  ), .I1 (nx34235z34
         ), .I2 (nx13298z15)) ;
         defparam ix12903z1706.INIT = 8'h96;
    LUT5 ix3326z39821 (.O (nx3326z3), .I0 (\plaintext(62)  ), .I1 (
         \p_key_samp(23)  ), .I2 (nx37232z13), .I3 (nx36230z11), .I4 (nx9305z10)
         ) ;
         defparam ix3326z39821.INIT = 32'h69969669;
    LUT6 ix9305z52044 (.O (nx9305z10), .I0 (nx13298z71), .I1 (nx13298z75), .I2 (
         nx13298z77), .I3 (nx13298z73), .I4 (nx13298z78), .I5 (nx13298z74)) ;
         defparam ix9305z52044.INIT = 64'h5267BCCB95CAC621;
    (* HLUTNM = "LUT62_1_65" *)
    LUT3 ix12903z1658 (.O (nx12903z258), .I0 (\plaintext(62)  ), .I1 (nx37232z13
         ), .I2 (nx36230z11)) ;
         defparam ix12903z1658.INIT = 8'h69;
    LUT5 ix3326z28345 (.O (nx3326z2), .I0 (\plaintext(30)  ), .I1 (
         \p_key_samp(38)  ), .I2 (nx63157z44), .I3 (px3752), .I4 (px3523)) ;
         defparam ix3326z28345.INIT = 32'h96696996;
    (* HLUTNM = "LUT62_1_43" *)
    LUT3 ix12903z1621 (.O (nx12903z214), .I0 (\plaintext(11)  ), .I1 (nx16286z6)
         , .I2 (nx13298z76)) ;
         defparam ix12903z1621.INIT = 8'h69;
    (* HLUTNM = "LUT62_1_4" *)
    LUT4 ix12903z28346 (.O (nx12903z3), .I0 (\plaintext(22)  ), .I1 (nx63157z4)
         , .I2 (nx37234z3), .I3 (nx11304z3)) ;
         defparam ix12903z28346.INIT = 16'h6996;
    (* HLUTNM = "LUT62_1_32" *)
    LUT4 ix22271z28344 (.O (px3503), .I0 (p_nbus_plaintext[63]), .I1 (nx63157z2)
         , .I2 (px3724), .I3 (px3504)) ;
         defparam ix22271z28344.INIT = 16'h6996;
    LUT6 ix22272z33160 (.O (px3504), .I0 (nx11304z2), .I1 (nx11304z4), .I2 (
         nx11304z5), .I3 (nx11304z7), .I4 (nx11304z8), .I5 (nx11304z9)) ;
         defparam ix22272z33160.INIT = 64'h37C78919C22D7C66;
    LUT5 ix11304z28352 (.O (nx11304z9), .I0 (plaintext[0]), .I1 (
         \p_key_samp(20)  ), .I2 (nx63157z28), .I3 (px3739), .I4 (px3506)) ;
         defparam ix11304z28352.INIT = 32'h96696996;
    LUT6 ix22274z55131 (.O (px3506), .I0 (nx7312z10), .I1 (nx7312z11), .I2 (
         nx7312z13), .I3 (nx7312z14), .I4 (nx7312z15), .I5 (nx7312z16)) ;
         defparam ix22274z55131.INIT = 64'h32D40D6B792ED239;
    LUT4 ix7312z39834 (.O (nx7312z16), .I0 (\plaintext(53)  ), .I1 (
         \p_key_samp(28)  ), .I2 (nx16289z10), .I3 (nx7312z17)) ;
         defparam ix7312z39834.INIT = 16'h9669;
    LUT6 ix7312z27559 (.O (nx7312z17), .I0 (nx24265z4), .I1 (nx24265z6), .I2 (
         nx24265z8), .I3 (nx24265z9), .I4 (nx24265z10), .I5 (nx24265z11)) ;
         defparam ix7312z27559.INIT = 64'h695946AABC866675;
    (* HLUTNM = "LUT62_1_96" *)
    LUT2 ix12903z2070 (.O (nx12903z429), .I0 (\plaintext(53)  ), .I1 (nx16289z10
         )) ;
         defparam ix12903z2070.INIT = 4'h9;
    LUT4 ix7312z28358 (.O (nx7312z15), .I0 (\plaintext(29)  ), .I1 (
         \p_key_samp(61)  ), .I2 (nx23267z2), .I3 (px3511)) ;
         defparam ix7312z28358.INIT = 16'h6996;
    LUT6 ix13298z50106 (.O (px3511), .I0 (nx24265z30), .I1 (nx24265z29), .I2 (
         nx24265z27), .I3 (nx24265z34), .I4 (nx24265z28), .I5 (nx24265z32)) ;
         defparam ix13298z50106.INIT = 64'h79B2864D600EBE79;
    (* HLUTNM = "LUT62_1_97" *)
    LUT2 ix23267z1320 (.O (px3512), .I0 (\plaintext(29)  ), .I1 (nx23267z2)) ;
         defparam ix23267z1320.INIT = 4'h6;
    LUT4 ix7312z39832 (.O (nx7312z14), .I0 (\p_plaintext(37)  ), .I1 (
         \p_key_samp(54)  ), .I2 (px3745), .I3 (px3514)) ;
         defparam ix7312z39832.INIT = 16'h9669;
    LUT6 ix13298z39551 (.O (px3514), .I0 (nx13298z12), .I1 (nx13298z14), .I2 (
         nx13298z16), .I3 (nx13298z17), .I4 (nx13298z18), .I5 (nx13298z19)) ;
         defparam ix13298z39551.INIT = 64'hC3966AC96A65953A;
    (* HLUTNM = "LUT62_1_97" *)
    LUT2 ix23270z1320 (.O (px3515), .I0 (\p_plaintext(37)  ), .I1 (px3745)) ;
         defparam ix23270z1320.INIT = 4'h6;
    LUT4 ix7312z39831 (.O (nx7312z13), .I0 (\plaintext(61)  ), .I1 (
         \p_key_samp(37)  ), .I2 (nx37232z2), .I3 (px3632)) ;
         defparam ix7312z39831.INIT = 16'h9669;
    LUT4 ix7312z28354 (.O (nx7312z11), .I0 (\plaintext(45)  ), .I1 (
         \p_key_samp(55)  ), .I2 (nx16289z7), .I3 (nx7312z12)) ;
         defparam ix7312z28354.INIT = 16'h6996;
    LUT6 ix7312z29379 (.O (nx7312z12), .I0 (nx24265z18), .I1 (nx24265z22), .I2 (
         nx24265z19), .I3 (nx24265z21), .I4 (nx24265z17), .I5 (nx24265z24)) ;
         defparam ix7312z29379.INIT = 64'hAD367289C2596D96;
    (* HLUTNM = "LUT62_1_90" *)
    LUT2 ix12903z1699 (.O (nx12903z435), .I0 (\plaintext(45)  ), .I1 (nx16289z7)
         ) ;
         defparam ix12903z1699.INIT = 4'h9;
    LUT4 ix7312z28353 (.O (nx7312z10), .I0 (plaintext[3]), .I1 (\p_key_samp(14)  
         ), .I2 (nx38222z2), .I3 (px3649)) ;
         defparam ix7312z28353.INIT = 16'h6996;
    (* HLUTNM = "LUT62_1_88" *)
    LUT3 ix24263z1464 (.O (px3521), .I0 (plaintext[0]), .I1 (nx63157z28), .I2 (
         px3739)) ;
         defparam ix24263z1464.INIT = 8'h96;
    LUT5 ix11304z28351 (.O (nx11304z8), .I0 (\plaintext(30)  ), .I1 (
         \p_key_samp(22)  ), .I2 (nx63157z44), .I3 (px3752), .I4 (px3523)) ;
         defparam ix11304z28351.INIT = 32'h96696996;
    LUT6 ix24265z13760 (.O (px3523), .I0 (nx24265z2), .I1 (nx24265z13), .I2 (
         nx24265z15), .I3 (nx24265z25), .I4 (nx24265z35), .I5 (nx24265z36)) ;
         defparam ix24265z13760.INIT = 64'h3C9ACBA5C9A5309E;
    LUT4 ix24265z28379 (.O (nx24265z36), .I0 (\plaintext(51)  ), .I1 (
         \p_key_samp(36)  ), .I2 (nx25263z8), .I3 (nx24265z37)) ;
         defparam ix24265z28379.INIT = 16'h6996;
    LUT6 ix24265z43025 (.O (nx24265z37), .I0 (nx37234z6), .I1 (nx37234z2), .I2 (
         nx37234z4), .I3 (nx37234z9), .I4 (nx37234z8), .I5 (nx37234z5)) ;
         defparam ix24265z43025.INIT = 64'h55E96935C316A2CB;
    (* HLUTNM = "LUT62_1_91" *)
    LUT2 ix12903z1703 (.O (nx12903z441), .I0 (\plaintext(51)  ), .I1 (nx25263z8)
         ) ;
         defparam ix12903z1703.INIT = 4'h6;
    LUT4 ix24265z39853 (.O (nx24265z35), .I0 (\plaintext(27)  ), .I1 (
         \p_key_samp(10)  ), .I2 (nx36228z2), .I3 (px3615)) ;
         defparam ix24265z39853.INIT = 16'h9669;
    LUT4 ix24265z28368 (.O (nx24265z25), .I0 (\plaintext(43)  ), .I1 (
         \p_key_samp(17)  ), .I2 (nx25263z6), .I3 (nx24265z26)) ;
         defparam ix24265z28368.INIT = 16'h6996;
    LUT6 ix24265z9212 (.O (nx24265z26), .I0 (nx24265z27), .I1 (nx24265z28), .I2 (
         nx24265z29), .I3 (nx24265z30), .I4 (nx24265z32), .I5 (nx24265z34)) ;
         defparam ix24265z9212.INIT = 64'hAA5A43B579A61EC1;
    (* HLUTNM = "LUT62_1_96" *)
    LUT2 ix12903z2095 (.O (nx12903z446), .I0 (\plaintext(43)  ), .I1 (nx25263z6)
         ) ;
         defparam ix12903z2095.INIT = 4'h6;
    LUT4 ix24265z39833 (.O (nx24265z15), .I0 (plaintext[5]), .I1 (
         \p_key_samp(60)  ), .I2 (nx27254z7), .I3 (px3543)) ;
         defparam ix24265z39833.INIT = 16'h9669;
    LUT4 ix24265z39831 (.O (nx24265z13), .I0 (\plaintext(59)  ), .I1 (
         \p_key_samp(34)  ), .I2 (nx27254z4), .I3 (px3546)) ;
         defparam ix24265z39831.INIT = 16'h9669;
    LUT4 ix24265z39820 (.O (nx24265z2), .I0 (\plaintext(35)  ), .I1 (
         \p_key_samp(27)  ), .I2 (nx39226z2), .I3 (px3652)) ;
         defparam ix24265z39820.INIT = 16'h9669;
    (* HLUTNM = "LUT62_1_89" *)
    LUT3 ix25263z1464 (.O (px3534), .I0 (\plaintext(30)  ), .I1 (nx63157z44), .I2 (
         px3752)) ;
         defparam ix25263z1464.INIT = 8'h96;
    LUT5 ix11304z28350 (.O (nx11304z7), .I0 (\plaintext(56)  ), .I1 (
         \p_key_samp(61)  ), .I2 (nx63157z20), .I3 (nx27254z2), .I4 (px3536)) ;
         defparam ix11304z28350.INIT = 32'h96696996;
    LUT6 ix25265z46896 (.O (px3536), .I0 (nx13298z4), .I1 (nx13298z6), .I2 (
         nx13298z7), .I3 (nx13298z8), .I4 (nx13298z10), .I5 (nx13298z20)) ;
         defparam ix25265z46896.INIT = 64'hB88767685E69B20E;
    LUT4 ix13298z28364 (.O (nx13298z20), .I0 (\plaintext(33)  ), .I1 (
         \p_key_samp(33)  ), .I2 (nx34235z10), .I3 (px3584)) ;
         defparam ix13298z28364.INIT = 16'h6996;
    LUT4 ix13298z28353 (.O (nx13298z10), .I0 (\plaintext(25)  ), .I1 (
         \p_key_samp(42)  ), .I2 (nx34235z31), .I3 (px3590)) ;
         defparam ix13298z28353.INIT = 16'h6996;
    LUT4 ix13298z28351 (.O (nx13298z8), .I0 (\plaintext(17)  ), .I1 (
         \p_key_samp(57)  ), .I2 (nx27254z11), .I3 (nx13298z9)) ;
         defparam ix13298z28351.INIT = 16'h6996;
    LUT6 ix13298z16907 (.O (nx13298z9), .I0 (nx24265z4), .I1 (nx24265z6), .I2 (
         nx24265z8), .I3 (nx24265z9), .I4 (nx24265z10), .I5 (nx24265z11)) ;
         defparam ix13298z16907.INIT = 64'h619E694B6A653CE1;
    (* HLUTNM = "LUT62_1_77" *)
    LUT2 ix12903z1586 (.O (nx12903z288), .I0 (\plaintext(17)  ), .I1 (nx27254z11
         )) ;
         defparam ix12903z1586.INIT = 4'h9;
    LUT4 ix13298z39825 (.O (nx13298z7), .I0 (plaintext[5]), .I1 (\p_key_samp(1)  
         ), .I2 (nx27254z7), .I3 (px3543)) ;
         defparam ix13298z39825.INIT = 16'h9669;
    LUT6 ix24265z8409 (.O (px3543), .I0 (nx24265z17), .I1 (nx24265z18), .I2 (
         nx24265z19), .I3 (nx24265z21), .I4 (nx24265z22), .I5 (nx24265z24)) ;
         defparam ix24265z8409.INIT = 64'hD3C3E44B6C171BA8;
    (* HLUTNM = "LUT62_1_98" *)
    LUT2 ix26260z1323 (.O (px3544), .I0 (plaintext[5]), .I1 (nx27254z7)) ;
         defparam ix26260z1323.INIT = 4'h9;
    LUT4 ix13298z39824 (.O (nx13298z6), .I0 (\plaintext(59)  ), .I1 (
         \p_key_samp(59)  ), .I2 (nx27254z4), .I3 (px3546)) ;
         defparam ix13298z39824.INIT = 16'h9669;
    LUT6 ix24265z12949 (.O (px3546), .I0 (nx36230z6), .I1 (nx36230z2), .I2 (
         nx36230z9), .I3 (nx36230z4), .I4 (nx36230z8), .I5 (nx36230z10)) ;
         defparam ix24265z12949.INIT = 64'h2CD3D22DD6A82D66;
    (* HLUTNM = "LUT62_1_98" *)
    LUT2 ix26263z1323 (.O (px3547), .I0 (\plaintext(59)  ), .I1 (nx27254z4)) ;
         defparam ix26263z1323.INIT = 4'h9;
    LUT4 ix13298z28347 (.O (nx13298z4), .I0 (\plaintext(9)  ), .I1 (
         \p_key_samp(19)  ), .I2 (nx27254z9), .I3 (nx13298z5)) ;
         defparam ix13298z28347.INIT = 16'h6996;
    LUT6 ix13298z41335 (.O (nx13298z5), .I0 (nx15291z3), .I1 (nx15291z13), .I2 (
         nx15291z15), .I3 (nx15291z25), .I4 (nx15291z35), .I5 (nx15291z37)) ;
         defparam ix13298z41335.INIT = 64'h69E7C63617A89C51;
    (* HLUTNM = "LUT62_1_74" *)
    LUT2 ix12903z1566 (.O (nx12903z265), .I0 (\plaintext(9)  ), .I1 (nx27254z9)
         ) ;
         defparam ix12903z1566.INIT = 4'h6;
    (* HLUTNM = "LUT62_1_90" *)
    LUT3 ix27254z1464 (.O (px3551), .I0 (\plaintext(56)  ), .I1 (nx63157z20), .I2 (
         nx27254z2)) ;
         defparam ix27254z1464.INIT = 8'h96;
    LUT5 ix11304z39823 (.O (nx11304z5), .I0 (\plaintext(14)  ), .I1 (
         \p_key_samp(37)  ), .I2 (nx63157z12), .I3 (nx37234z7), .I4 (nx11304z6)
         ) ;
         defparam ix11304z39823.INIT = 32'h69969669;
    LUT6 ix11304z35856 (.O (nx11304z6), .I0 (nx13298z38), .I1 (nx13298z40), .I2 (
         nx13298z41), .I3 (nx13298z42), .I4 (nx13298z44), .I5 (nx13298z45)) ;
         defparam ix11304z35856.INIT = 64'h23DDE817782986E9;
    LUT4 ix13298z28389 (.O (nx13298z45), .I0 (\plaintext(47)  ), .I1 (
         \p_key_samp(53)  ), .I2 (nx15291z12), .I3 (nx13298z46)) ;
         defparam ix13298z28389.INIT = 16'h6996;
    LUT6 ix13298z43660 (.O (nx13298z46), .I0 (nx36230z2), .I1 (nx36230z4), .I2 (
         nx36230z6), .I3 (nx36230z8), .I4 (nx36230z9), .I5 (nx36230z10)) ;
         defparam ix13298z43660.INIT = 64'hB51A69365AC3A53C;
    (* HLUTNM = "LUT62_1_89" *)
    LUT2 ix12903z1679 (.O (nx12903z410), .I0 (\plaintext(47)  ), .I1 (nx15291z12
         )) ;
         defparam ix12903z1679.INIT = 4'h6;
    LUT4 ix13298z39863 (.O (nx13298z44), .I0 (p_nbus_plaintext[63]), .I1 (
         \p_key_samp(13)  ), .I2 (nx63157z2), .I3 (px3724)) ;
         defparam ix13298z39863.INIT = 16'h9669;
    LUT4 ix13298z28386 (.O (nx13298z42), .I0 (\p_plaintext(39)  ), .I1 (
         \p_key_samp(63)  ), .I2 (px3781), .I3 (px3559)) ;
         defparam ix13298z28386.INIT = 16'h6996;
    LUT6 ix13298z57268 (.O (px3559), .I0 (nx24265z4), .I1 (nx24265z6), .I2 (
         nx24265z8), .I3 (nx24265z9), .I4 (nx24265z10), .I5 (nx24265z11)) ;
         defparam ix13298z57268.INIT = 64'hD947219C29E8DA67;
    (* HLUTNM = "LUT62_1_99" *)
    LUT2 ix28250z1320 (.O (px3560), .I0 (\p_plaintext(39)  ), .I1 (px3781)) ;
         defparam ix28250z1320.INIT = 4'h6;
    LUT4 ix13298z28385 (.O (nx13298z41), .I0 (\plaintext(31)  ), .I1 (
         \p_key_samp(22)  ), .I2 (nx28253z2), .I3 (px3562)) ;
         defparam ix13298z28385.INIT = 16'h6996;
    LUT6 ix7313z15849 (.O (px3562), .I0 (nx7313z3), .I1 (nx7313z5), .I2 (
         nx7313z6), .I3 (nx7313z8), .I4 (nx7313z9), .I5 (nx7313z11)) ;
         defparam ix7313z15849.INIT = 64'h97466D9BC23538C6;
    (* HLUTNM = "LUT62_1_99" *)
    LUT2 ix28253z1320 (.O (px3563), .I0 (\plaintext(31)  ), .I1 (nx28253z2)) ;
         defparam ix28253z1320.INIT = 4'h6;
    LUT4 ix13298z39859 (.O (nx13298z40), .I0 (\p_plaintext(63)  ), .I1 (
         \p_key_samp(7)  ), .I2 (nx29253z2), .I3 (px3565)) ;
         defparam ix13298z39859.INIT = 16'h9669;
    LUT6 ix13298z31496 (.O (px3565), .I0 (nx24265z17), .I1 (nx24265z19), .I2 (
         nx24265z18), .I3 (nx24265z22), .I4 (nx24265z21), .I5 (nx24265z24)) ;
         defparam ix13298z31496.INIT = 64'hC16E9A8716B075CB;
    LUT4 ix24265z28367 (.O (nx24265z24), .I0 (plaintext[4]), .I1 (
         \p_key_samp(9)  ), .I2 (nx36228z6), .I3 (px3626)) ;
         defparam ix24265z28367.INIT = 16'h6996;
    LUT4 ix24265z28364 (.O (nx24265z21), .I0 (\plaintext(26)  ), .I1 (
         \p_key_samp(36)  ), .I2 (nx45210z2), .I3 (px3716)) ;
         defparam ix24265z28364.INIT = 16'h6996;
    LUT4 ix24265z39840 (.O (nx24265z22), .I0 (\plaintext(10)  ), .I1 (
         \p_key_samp(2)  ), .I2 (nx29253z10), .I3 (nx24265z23)) ;
         defparam ix24265z39840.INIT = 16'h9669;
    LUT6 ix24265z36660 (.O (nx24265z23), .I0 (nx15291z5), .I1 (nx15291z6), .I2 (
         nx15291z7), .I3 (nx15291z9), .I4 (nx15291z10), .I5 (nx15291z11)) ;
         defparam ix24265z36660.INIT = 64'hD29E6712871689FC;
    (* HLUTNM = "LUT62_1_73" *)
    LUT2 ix12903z1548 (.O (nx12903z241), .I0 (\plaintext(10)  ), .I1 (nx29253z10
         )) ;
         defparam ix12903z1548.INIT = 4'h9;
    LUT4 ix24265z39836 (.O (nx24265z18), .I0 (\plaintext(60)  ), .I1 (
         \p_key_samp(19)  ), .I2 (nx36228z10), .I3 (px3623)) ;
         defparam ix24265z39836.INIT = 16'h9669;
    LUT4 ix24265z39837 (.O (nx24265z19), .I0 (\plaintext(18)  ), .I1 (
         \p_key_samp(50)  ), .I2 (nx29253z8), .I3 (nx24265z20)) ;
         defparam ix24265z39837.INIT = 16'h9669;
    LUT6 ix24265z22779 (.O (nx24265z20), .I0 (nx25263z3), .I1 (nx25263z4), .I2 (
         nx25263z5), .I3 (nx25263z7), .I4 (nx25263z9), .I5 (nx25263z10)) ;
         defparam ix24265z22779.INIT = 64'hA9746C39A96353C6;
    (* HLUTNM = "LUT62_1_92" *)
    LUT2 ix12903z1747 (.O (nx12903z227), .I0 (\plaintext(18)  ), .I1 (nx29253z8)
         ) ;
         defparam ix12903z1747.INIT = 4'h6;
    LUT4 ix24265z28360 (.O (nx24265z17), .I0 (\plaintext(34)  ), .I1 (
         \p_key_samp(33)  ), .I2 (nx41222z2), .I3 (px3688)) ;
         defparam ix24265z28360.INIT = 16'h6996;
    (* HLUTNM = "LUT62_1_100" *)
    LUT2 ix29253z1323 (.O (px3576), .I0 (\p_plaintext(63)  ), .I1 (nx29253z2)) ;
         defparam ix29253z1323.INIT = 4'h9;
    LUT4 ix13298z28382 (.O (nx13298z38), .I0 (\plaintext(55)  ), .I1 (
         \p_key_samp(46)  ), .I2 (nx15291z8), .I3 (nx13298z39)) ;
         defparam ix13298z28382.INIT = 16'h6996;
    LUT6 ix13298z13098 (.O (nx13298z39), .I0 (nx24265z27), .I1 (nx24265z30), .I2 (
         nx24265z29), .I3 (nx24265z28), .I4 (nx24265z34), .I5 (nx24265z32)) ;
         defparam ix13298z13098.INIT = 64'h3D92D22D926B2DE1;
    (* HLUTNM = "LUT62_1_87" *)
    LUT2 ix12903z1670 (.O (nx12903z395), .I0 (\plaintext(55)  ), .I1 (nx15291z8)
         ) ;
         defparam ix12903z1670.INIT = 4'h9;
    (* HLUTNM = "LUT62_1_95" *)
    LUT3 ix61487z1468 (.O (nx61487z6), .I0 (\plaintext(14)  ), .I1 (nx63157z12)
         , .I2 (nx37234z7)) ;
         defparam ix61487z1468.INIT = 8'h96;
    LUT5 ix11304z28347 (.O (nx11304z4), .I0 (\plaintext(38)  ), .I1 (
         \p_key_samp(54)  ), .I2 (nx63157z36), .I3 (px3726), .I4 (px3582)) ;
         defparam ix11304z28347.INIT = 32'h96696996;
    LUT6 ix30246z15209 (.O (px3582), .I0 (nx13298z61), .I1 (nx13298z63), .I2 (
         nx13298z64), .I3 (nx13298z66), .I4 (nx13298z67), .I5 (nx13298z68)) ;
         defparam ix30246z15209.INIT = 64'h9678D2A9E12E3647;
    LUT4 ix13298z28412 (.O (nx13298z68), .I0 (\plaintext(33)  ), .I1 (
         \p_key_samp(43)  ), .I2 (nx34235z10), .I3 (px3584)) ;
         defparam ix13298z28412.INIT = 16'h6996;
    LUT6 ix13298z58965 (.O (px3584), .I0 (nx7313z11), .I1 (nx7313z9), .I2 (
         nx7313z3), .I3 (nx7313z8), .I4 (nx7313z6), .I5 (nx7313z5)) ;
         defparam ix13298z58965.INIT = 64'hA59E4E612E59E11E;
    (* HLUTNM = "LUT62_1_100" *)
    LUT2 ix30249z1320 (.O (px3585), .I0 (\plaintext(33)  ), .I1 (nx34235z10)) ;
         defparam ix30249z1320.INIT = 4'h6;
    LUT4 ix13298z28411 (.O (nx13298z67), .I0 (\plaintext(7)  ), .I1 (
         \p_key_samp(26)  ), .I2 (nx34235z6), .I3 (px3587)) ;
         defparam ix13298z28411.INIT = 16'h6996;
    LUT6 ix13298z57539 (.O (px3587), .I0 (nx15291z3), .I1 (nx15291z13), .I2 (
         nx15291z15), .I3 (nx15291z25), .I4 (nx15291z35), .I5 (nx15291z37)) ;
         defparam ix13298z57539.INIT = 64'h45362AD49C93DB69;
    (* HLUTNM = "LUT62_1_101" *)
    LUT2 ix30252z1320 (.O (px3588), .I0 (\plaintext(7)  ), .I1 (nx34235z6)) ;
         defparam ix30252z1320.INIT = 4'h6;
    LUT4 ix13298z28410 (.O (nx13298z66), .I0 (\plaintext(25)  ), .I1 (
         \p_key_samp(44)  ), .I2 (nx34235z31), .I3 (px3590)) ;
         defparam ix13298z28410.INIT = 16'h6996;
    LUT6 ix13298z22744 (.O (px3590), .I0 (nx13298z12), .I1 (nx13298z14), .I2 (
         nx13298z16), .I3 (nx13298z17), .I4 (nx13298z18), .I5 (nx13298z19)) ;
         defparam ix13298z22744.INIT = 64'h4EB13C5339C653AC;
    (* HLUTNM = "LUT62_1_101" *)
    LUT2 ix31242z1320 (.O (px3591), .I0 (\plaintext(25)  ), .I1 (nx34235z31)) ;
         defparam ix31242z1320.INIT = 4'h6;
    LUT4 ix13298z39883 (.O (nx13298z64), .I0 (\plaintext(41)  ), .I1 (
         \p_key_samp(9)  ), .I2 (nx34235z8), .I3 (nx13298z65)) ;
         defparam ix13298z39883.INIT = 16'h9669;
    LUT6 ix13298z36538 (.O (nx13298z65), .I0 (nx36230z2), .I1 (nx36230z4), .I2 (
         nx36230z6), .I3 (nx36230z8), .I4 (nx36230z9), .I5 (nx36230z10)) ;
         defparam ix13298z36538.INIT = 64'hA6D153E496658957;
    (* HLUTNM = "LUT62_1_85" *)
    LUT2 ix12903z1631 (.O (nx12903z347), .I0 (\plaintext(41)  ), .I1 (nx34235z8)
         ) ;
         defparam ix12903z1631.INIT = 4'h9;
    LUT4 ix13298z28407 (.O (nx13298z63), .I0 (\plaintext(57)  ), .I1 (
         \p_key_samp(2)  ), .I2 (nx34235z21), .I3 (px3596)) ;
         defparam ix13298z28407.INIT = 16'h6996;
    LUT6 ix13298z13036 (.O (px3596), .I0 (nx24265z30), .I1 (nx24265z29), .I2 (
         nx24265z27), .I3 (nx24265z34), .I4 (nx24265z28), .I5 (nx24265z32)) ;
         defparam ix13298z13036.INIT = 64'h9DE8E25B920B2D96;
    LUT4 ix24265z28375 (.O (nx24265z32), .I0 (\plaintext(16)  ), .I1 (
         \p_key_samp(41)  ), .I2 (nx34235z28), .I3 (nx24265z33)) ;
         defparam ix24265z28375.INIT = 16'h6996;
    LUT6 ix24265z27563 (.O (nx24265z33), .I0 (nx34235z3), .I1 (nx34235z5), .I2 (
         nx34235z7), .I3 (nx34235z9), .I4 (nx34235z20), .I5 (nx34235z30)) ;
         defparam ix24265z27563.INIT = 64'h788647B93C996669;
    (* HLUTNM = "LUT62_1_88" *)
    LUT2 ix12903z1678 (.O (nx12903z404), .I0 (\plaintext(16)  ), .I1 (nx34235z28
         )) ;
         defparam ix12903z1678.INIT = 4'h9;
    LUT4 ix24265z28371 (.O (nx24265z28), .I0 (\plaintext(24)  ), .I1 (
         \p_key_samp(26)  ), .I2 (nx39226z17), .I3 (px3657)) ;
         defparam ix24265z28371.INIT = 16'h6996;
    LUT4 ix24265z28377 (.O (nx24265z34), .I0 (\plaintext(32)  ), .I1 (
         \p_key_samp(17)  ), .I2 (nx39226z15), .I3 (px3665)) ;
         defparam ix24265z28377.INIT = 16'h6996;
    LUT4 ix24265z39845 (.O (nx24265z27), .I0 (plaintext[6]), .I1 (
         \p_key_samp(52)  ), .I2 (nx44209z2), .I3 (px3702)) ;
         defparam ix24265z39845.INIT = 16'h9669;
    LUT4 ix24265z28372 (.O (nx24265z29), .I0 (\plaintext(58)  ), .I1 (
         \p_key_samp(43)  ), .I2 (nx34235z18), .I3 (px3705)) ;
         defparam ix24265z28372.INIT = 16'h6996;
    LUT4 ix24265z28373 (.O (nx24265z30), .I0 (\plaintext(8)  ), .I1 (
         \p_key_samp(3)  ), .I2 (nx34235z25), .I3 (nx24265z31)) ;
         defparam ix24265z28373.INIT = 16'h6996;
    LUT6 ix24265z52691 (.O (nx24265z31), .I0 (nx16289z4), .I1 (nx16289z8), .I2 (
         nx16289z3), .I3 (px3744), .I4 (nx16289z6), .I5 (nx16289z9)) ;
         defparam ix24265z52691.INIT = 64'h1EB4790CA779C893;
    (* HLUTNM = "LUT62_1_95" *)
    LUT2 ix12903z2023 (.O (nx12903z400), .I0 (\plaintext(8)  ), .I1 (nx34235z25)
         ) ;
         defparam ix12903z2023.INIT = 4'h6;
    (* HLUTNM = "LUT62_1_102" *)
    LUT2 ix33244z1320 (.O (px3607), .I0 (\plaintext(57)  ), .I1 (nx34235z21)) ;
         defparam ix33244z1320.INIT = 4'h6;
    LUT4 ix13298z28405 (.O (nx13298z61), .I0 (\plaintext(49)  ), .I1 (
         \p_key_samp(58)  ), .I2 (nx34235z4), .I3 (nx13298z62)) ;
         defparam ix13298z28405.INIT = 16'h6996;
    LUT6 ix13298z28413 (.O (nx13298z62), .I0 (nx37234z2), .I1 (nx37234z4), .I2 (
         nx37234z6), .I3 (nx37234z9), .I4 (nx37234z5), .I5 (nx37234z8)) ;
         defparam ix13298z28413.INIT = 64'h69C31E59C722699D;
    (* HLUTNM = "LUT62_1_82" *)
    LUT2 ix12903z1619 (.O (nx12903z335), .I0 (\plaintext(49)  ), .I1 (nx34235z4)
         ) ;
         defparam ix12903z1619.INIT = 4'h6;
    (* HLUTNM = "LUT62_1_91" *)
    LUT3 ix34235z1464 (.O (px3611), .I0 (\plaintext(38)  ), .I1 (nx63157z36), .I2 (
         px3726)) ;
         defparam ix34235z1464.INIT = 8'h96;
    LUT5 ix11304z28345 (.O (nx11304z2), .I0 (\plaintext(22)  ), .I1 (
         \p_key_samp(47)  ), .I2 (nx63157z4), .I3 (nx37234z3), .I4 (nx11304z3)
         ) ;
         defparam ix11304z28345.INIT = 32'h96696996;
    LUT6 ix11304z19837 (.O (nx11304z3), .I0 (nx13298z71), .I1 (nx13298z75), .I2 (
         nx13298z77), .I3 (nx13298z73), .I4 (nx13298z78), .I5 (nx13298z74)) ;
         defparam ix11304z19837.INIT = 64'h89737EA5B42D4859;
    LUT4 ix13298z39893 (.O (nx13298z74), .I0 (\plaintext(27)  ), .I1 (
         \p_key_samp(52)  ), .I2 (nx36228z2), .I3 (px3615)) ;
         defparam ix13298z39893.INIT = 16'h9669;
    LUT6 ix15291z16136 (.O (px3615), .I0 (nx15291z3), .I1 (nx15291z13), .I2 (
         nx15291z15), .I3 (nx15291z25), .I4 (nx15291z35), .I5 (nx15291z37)) ;
         defparam ix15291z16136.INIT = 64'h668E9C93817A39E5;
    LUT4 ix15291z28379 (.O (nx15291z37), .I0 (\plaintext(44)  ), .I1 (
         \p_key_samp(39)  ), .I2 (nx36228z4), .I3 (nx15291z38)) ;
         defparam ix15291z28379.INIT = 16'h6996;
    LUT6 ix15291z46771 (.O (nx15291z38), .I0 (nx16286z8), .I1 (nx16286z7), .I2 (
         nx16286z3), .I3 (nx16286z5), .I4 (nx16286z10), .I5 (nx16286z4)) ;
         defparam ix15291z46771.INIT = 64'h923D5E866C92B16D;
    (* HLUTNM = "LUT62_1_76" *)
    LUT2 ix12903z1583 (.O (nx12903z283), .I0 (\plaintext(44)  ), .I1 (nx36228z4)
         ) ;
         defparam ix12903z1583.INIT = 4'h9;
    LUT4 ix15291z28377 (.O (nx15291z35), .I0 (\plaintext(52)  ), .I1 (
         \p_key_samp(12)  ), .I2 (nx36228z8), .I3 (nx15291z36)) ;
         defparam ix15291z28377.INIT = 16'h6996;
    LUT6 ix15291z25326 (.O (nx15291z36), .I0 (nx34235z3), .I1 (nx34235z5), .I2 (
         nx34235z7), .I3 (nx34235z9), .I4 (nx34235z20), .I5 (nx34235z30)) ;
         defparam ix15291z25326.INIT = 64'h9EE12669700F5DAA;
    (* HLUTNM = "LUT62_1_75" *)
    LUT2 ix12903z1572 (.O (nx12903z270), .I0 (\plaintext(52)  ), .I1 (nx36228z8)
         ) ;
         defparam ix12903z1572.INIT = 4'h9;
    LUT4 ix15291z39842 (.O (nx15291z25), .I0 (\plaintext(60)  ), .I1 (
         \p_key_samp(21)  ), .I2 (nx36228z10), .I3 (px3623)) ;
         defparam ix15291z39842.INIT = 16'h9669;
    LUT6 ix15291z22751 (.O (px3623), .I0 (nx15291z27), .I1 (nx15291z28), .I2 (
         nx15291z30), .I3 (nx15291z31), .I4 (nx15291z33), .I5 (nx15291z34)) ;
         defparam ix15291z22751.INIT = 64'h91B68D5A6C6953A5;
    (* HLUTNM = "LUT62_1_102" *)
    LUT2 ix35235z1323 (.O (px3624), .I0 (\plaintext(60)  ), .I1 (nx36228z10)) ;
         defparam ix35235z1323.INIT = 4'h9;
    LUT4 ix15291z28358 (.O (nx15291z15), .I0 (plaintext[4]), .I1 (
         \p_key_samp(63)  ), .I2 (nx36228z6), .I3 (px3626)) ;
         defparam ix15291z28358.INIT = 16'h6996;
    LUT6 ix15291z8876 (.O (px3626), .I0 (nx15291z17), .I1 (px3697), .I2 (
         nx15291z20), .I3 (nx15291z21), .I4 (nx15291z22), .I5 (nx15291z23)) ;
         defparam ix15291z8876.INIT = 64'hE53D90465AC11D7B;
    (* HLUTNM = "LUT62_1_103" *)
    LUT2 ix35238z1320 (.O (px3627), .I0 (plaintext[4]), .I1 (nx36228z6)) ;
         defparam ix35238z1320.INIT = 4'h6;
    LUT4 ix15291z39831 (.O (nx15291z13), .I0 (\plaintext(28)  ), .I1 (
         \p_key_samp(45)  ), .I2 (nx37232z9), .I3 (px3638)) ;
         defparam ix15291z39831.INIT = 16'h9669;
    LUT4 ix15291z39821 (.O (nx15291z3), .I0 (\plaintext(36)  ), .I1 (
         \p_key_samp(38)  ), .I2 (nx37232z11), .I3 (px3635)) ;
         defparam ix15291z39821.INIT = 16'h9669;
    (* HLUTNM = "LUT62_1_103" *)
    LUT2 ix36228z1323 (.O (px3630), .I0 (\plaintext(27)  ), .I1 (nx36228z2)) ;
         defparam ix36228z1323.INIT = 4'h9;
    LUT4 ix13298z39897 (.O (nx13298z78), .I0 (\plaintext(61)  ), .I1 (
         \p_key_samp(35)  ), .I2 (nx37232z2), .I3 (px3632)) ;
         defparam ix13298z39897.INIT = 16'h9669;
    LUT6 ix36230z18588 (.O (px3632), .I0 (nx36230z2), .I1 (nx36230z4), .I2 (
         nx36230z6), .I3 (nx36230z8), .I4 (nx36230z9), .I5 (nx36230z10)) ;
         defparam ix36230z18588.INIT = 64'h8B563CA57C29437A;
    LUT4 ix36230z39828 (.O (nx36230z10), .I0 (\plaintext(62)  ), .I1 (
         \p_key_samp(7)  ), .I2 (nx37232z13), .I3 (nx36230z11)) ;
         defparam ix36230z39828.INIT = 16'h9669;
    LUT4 ix36230z39827 (.O (nx36230z9), .I0 (\plaintext(36)  ), .I1 (
         \p_key_samp(46)  ), .I2 (nx37232z11), .I3 (px3635)) ;
         defparam ix36230z39827.INIT = 16'h9669;
    LUT6 ix15291z12958 (.O (px3635), .I0 (nx15291z5), .I1 (nx15291z6), .I2 (
         nx15291z7), .I3 (nx15291z9), .I4 (nx15291z10), .I5 (nx15291z11)) ;
         defparam ix15291z12958.INIT = 64'h6A59962CD1A62D79;
    (* HLUTNM = "LUT62_1_104" *)
    LUT2 ix36234z1320 (.O (px3636), .I0 (\plaintext(36)  ), .I1 (nx37232z11)) ;
         defparam ix36234z1320.INIT = 4'h6;
    LUT4 ix36230z39826 (.O (nx36230z8), .I0 (\plaintext(28)  ), .I1 (
         \p_key_samp(31)  ), .I2 (nx37232z9), .I3 (px3638)) ;
         defparam ix36230z39826.INIT = 16'h9669;
    LUT6 ix15291z39328 (.O (px3638), .I0 (nx27254z3), .I1 (nx27254z5), .I2 (
         nx27254z6), .I3 (nx27254z8), .I4 (nx27254z10), .I5 (nx27254z12)) ;
         defparam ix15291z39328.INIT = 64'h38146B8EDE6B9471;
    (* HLUTNM = "LUT62_1_104" *)
    LUT2 ix36237z1323 (.O (px3639), .I0 (\plaintext(28)  ), .I1 (nx37232z9)) ;
         defparam ix36237z1323.INIT = 4'h9;
    LUT4 ix36230z39824 (.O (nx36230z6), .I0 (plaintext[2]), .I1 (\p_key_samp(4)  
         ), .I2 (nx40221z2), .I3 (px3674)) ;
         defparam ix36230z39824.INIT = 16'h9669;
    LUT4 ix36230z28347 (.O (nx36230z4), .I0 (\plaintext(20)  ), .I1 (
         \p_key_samp(14)  ), .I2 (nx37232z6), .I3 (nx36230z5)) ;
         defparam ix36230z28347.INIT = 16'h6996;
    LUT6 ix36230z38803 (.O (nx36230z5), .I0 (nx25263z3), .I1 (nx25263z4), .I2 (
         nx25263z5), .I3 (nx25263z7), .I4 (nx25263z9), .I5 (nx25263z10)) ;
         defparam ix36230z38803.INIT = 64'hB658D8630DB6926D;
    (* HLUTNM = "LUT62_1_94" *)
    LUT2 ix12903z1945 (.O (nx12903z351), .I0 (\plaintext(20)  ), .I1 (nx37232z6)
         ) ;
         defparam ix12903z1945.INIT = 4'h6;
    LUT4 ix36230z39820 (.O (nx36230z2), .I0 (\plaintext(12)  ), .I1 (
         \p_key_samp(13)  ), .I2 (nx37232z4), .I3 (nx36230z3)) ;
         defparam ix36230z39820.INIT = 16'h9669;
    LUT6 ix36230z9176 (.O (nx36230z3), .I0 (nx16289z4), .I1 (nx16289z8), .I2 (
         nx16289z3), .I3 (px3744), .I4 (nx16289z6), .I5 (nx16289z9)) ;
         defparam ix36230z9176.INIT = 64'h896C70C7C79A1EB4;
    (* HLUTNM = "LUT62_1_86" *)
    LUT2 ix12903z1635 (.O (nx12903z355), .I0 (\plaintext(12)  ), .I1 (nx37232z4)
         ) ;
         defparam ix12903z1635.INIT = 4'h6;
    (* HLUTNM = "LUT62_1_105" *)
    LUT2 ix37232z1320 (.O (px3647), .I0 (\plaintext(61)  ), .I1 (nx37232z2)) ;
         defparam ix37232z1320.INIT = 4'h6;
    LUT4 ix13298z28417 (.O (nx13298z73), .I0 (plaintext[3]), .I1 (
         \p_key_samp(25)  ), .I2 (nx38222z2), .I3 (px3649)) ;
         defparam ix13298z28417.INIT = 16'h6996;
    LUT6 ix37234z28850 (.O (px3649), .I0 (nx37234z2), .I1 (nx37234z4), .I2 (
         nx37234z5), .I3 (nx37234z6), .I4 (nx37234z8), .I5 (nx37234z9)) ;
         defparam ix37234z28850.INIT = 64'h6768DA1E78996B90;
    (* HLUTNM = "LUT62_1_105" *)
    LUT2 ix38222z1320 (.O (px3650), .I0 (plaintext[3]), .I1 (nx38222z2)) ;
         defparam ix38222z1320.INIT = 4'h6;
    LUT4 ix13298z39896 (.O (nx13298z77), .I0 (\plaintext(35)  ), .I1 (
         \p_key_samp(49)  ), .I2 (nx39226z2), .I3 (px3652)) ;
         defparam ix13298z39896.INIT = 16'h9669;
    LUT6 ix24265z21194 (.O (px3652), .I0 (nx24265z4), .I1 (nx24265z6), .I2 (
         nx24265z8), .I3 (nx24265z9), .I4 (nx24265z10), .I5 (nx24265z11)) ;
         defparam ix24265z21194.INIT = 64'h1DD4E239A25E4DA6;
    LUT4 ix24265z39829 (.O (nx24265z11), .I0 (\plaintext(40)  ), .I1 (
         \p_key_samp(60)  ), .I2 (nx39226z7), .I3 (nx24265z12)) ;
         defparam ix24265z39829.INIT = 16'h9669;
    LUT6 ix24265z44165 (.O (nx24265z12), .I0 (nx15291z27), .I1 (nx15291z34), .I2 (
         nx15291z31), .I3 (nx15291z28), .I4 (nx15291z30), .I5 (nx15291z33)) ;
         defparam ix24265z44165.INIT = 64'h03D918D7D83EA758;
    (* HLUTNM = "LUT62_1_79" *)
    LUT2 ix12903z1593 (.O (nx12903z299), .I0 (\plaintext(40)  ), .I1 (nx39226z7)
         ) ;
         defparam ix12903z1593.INIT = 4'h6;
    LUT4 ix24265z28353 (.O (nx24265z10), .I0 (\plaintext(24)  ), .I1 (
         \p_key_samp(59)  ), .I2 (nx39226z17), .I3 (px3657)) ;
         defparam ix24265z28353.INIT = 16'h6996;
    LUT6 ix12297z40326 (.O (px3657), .I0 (nx15291z5), .I1 (nx15291z6), .I2 (
         nx15291z7), .I3 (nx15291z9), .I4 (nx15291z10), .I5 (nx15291z11)) ;
         defparam ix12297z40326.INIT = 64'h0BF4F44B6D929863;
    (* HLUTNM = "LUT62_1_106" *)
    LUT2 ix38230z1323 (.O (px3658), .I0 (\plaintext(24)  ), .I1 (nx39226z17)) ;
         defparam ix38230z1323.INIT = 4'h9;
    LUT4 ix24265z28352 (.O (nx24265z9), .I0 (\plaintext(56)  ), .I1 (
         \p_key_samp(49)  ), .I2 (nx63157z20), .I3 (nx27254z2)) ;
         defparam ix24265z28352.INIT = 16'h6996;
    LUT4 ix24265z28351 (.O (nx24265z8), .I0 (plaintext[0]), .I1 (
         \p_key_samp(10)  ), .I2 (nx63157z28), .I3 (px3739)) ;
         defparam ix24265z28351.INIT = 16'h6996;
    LUT4 ix24265z28349 (.O (nx24265z6), .I0 (\plaintext(48)  ), .I1 (
         \p_key_samp(42)  ), .I2 (nx39226z4), .I3 (nx24265z7)) ;
         defparam ix24265z28349.INIT = 16'h6996;
    LUT6 ix24265z59566 (.O (nx24265z7), .I0 (nx15291z22), .I1 (nx15291z21), .I2 (
         px3697), .I3 (nx15291z23), .I4 (nx15291z17), .I5 (nx15291z20)) ;
         defparam ix24265z59566.INIT = 64'hE79A54291675E386;
    (* HLUTNM = "LUT62_1_93" *)
    LUT2 ix12903z1855 (.O (nx12903z293), .I0 (\plaintext(48)  ), .I1 (nx39226z4)
         ) ;
         defparam ix12903z1855.INIT = 4'h6;
    LUT4 ix24265z28347 (.O (nx24265z4), .I0 (\plaintext(32)  ), .I1 (
         \p_key_samp(27)  ), .I2 (nx39226z15), .I3 (px3665)) ;
         defparam ix24265z28347.INIT = 16'h6996;
    LUT6 ix24265z47506 (.O (px3665), .I0 (nx25263z7), .I1 (nx25263z5), .I2 (
         nx25263z10), .I3 (nx25263z9), .I4 (nx25263z4), .I5 (nx25263z3)) ;
         defparam ix24265z47506.INIT = 64'hC32C69954ED3B46C;
    (* HLUTNM = "LUT62_1_106" *)
    LUT2 ix39225z1320 (.O (px3666), .I0 (\plaintext(32)  ), .I1 (nx39226z15)) ;
         defparam ix39225z1320.INIT = 4'h6;
    (* HLUTNM = "LUT62_1_107" *)
    LUT2 ix39226z1320 (.O (px3667), .I0 (\plaintext(35)  ), .I1 (nx39226z2)) ;
         defparam ix39226z1320.INIT = 4'h6;
    LUT4 ix13298z39894 (.O (nx13298z75), .I0 (\plaintext(11)  ), .I1 (
         \p_key_samp(18)  ), .I2 (nx16286z6), .I3 (nx13298z76)) ;
         defparam ix13298z39894.INIT = 16'h9669;
    LUT6 ix13298z16852 (.O (nx13298z76), .I0 (nx13298z12), .I1 (nx13298z14), .I2 (
         nx13298z16), .I3 (nx13298z17), .I4 (nx13298z18), .I5 (nx13298z19)) ;
         defparam ix13298z16852.INIT = 64'h595A5CA3A3C33C66;
    LUT4 ix13298z39838 (.O (nx13298z19), .I0 (\plaintext(62)  ), .I1 (
         \p_key_samp(20)  ), .I2 (nx37232z13), .I3 (nx36230z11)) ;
         defparam ix13298z39838.INIT = 16'h9669;
    LUT6 ix36230z15492 (.O (nx36230z11), .I0 (nx16286z4), .I1 (nx16286z7), .I2 (
         nx16286z8), .I3 (nx16286z3), .I4 (nx16286z5), .I5 (nx16286z10)) ;
         defparam ix36230z15492.INIT = 64'h2A95C1C69EE33758;
    (* HLUTNM = "LUT62_1_65" *)
    LUT2 ix12903z1482 (.O (nx12903z165), .I0 (\plaintext(62)  ), .I1 (nx37232z13
         )) ;
         defparam ix12903z1482.INIT = 4'h6;
    LUT4 ix13298z39856 (.O (nx13298z18), .I0 (plaintext[2]), .I1 (
         \p_key_samp(62)  ), .I2 (nx40221z2), .I3 (px3674)) ;
         defparam ix13298z39856.INIT = 16'h9669;
    LUT6 ix36230z17372 (.O (px3674), .I0 (nx15291z20), .I1 (nx15291z23), .I2 (
         px3697), .I3 (nx15291z17), .I4 (nx15291z22), .I5 (nx15291z21)) ;
         defparam ix36230z17372.INIT = 64'h5A3FA45981C33EB4;
    (* HLUTNM = "LUT62_1_107" *)
    LUT2 ix40221z1320 (.O (px3675), .I0 (plaintext[2]), .I1 (nx40221z2)) ;
         defparam ix40221z1320.INIT = 4'h6;
    LUT4 ix13298z28360 (.O (nx13298z17), .I0 (\plaintext(30)  ), .I1 (
         \p_key_samp(6)  ), .I2 (nx63157z44), .I3 (px3752)) ;
         defparam ix13298z28360.INIT = 16'h6996;
    LUT4 ix13298z28359 (.O (nx13298z16), .I0 (\plaintext(38)  ), .I1 (
         \p_key_samp(47)  ), .I2 (nx63157z36), .I3 (px3726)) ;
         defparam ix13298z28359.INIT = 16'h6996;
    LUT4 ix13298z28357 (.O (nx13298z14), .I0 (\plaintext(54)  ), .I1 (
         \p_key_samp(30)  ), .I2 (nx34235z34), .I3 (nx13298z15)) ;
         defparam ix13298z28357.INIT = 16'h6996;
    LUT6 ix13298z41105 (.O (nx13298z15), .I0 (nx27254z8), .I1 (nx27254z6), .I2 (
         nx27254z5), .I3 (nx27254z10), .I4 (nx27254z12), .I5 (nx27254z3)) ;
         defparam ix13298z41105.INIT = 64'h1EE1741E615E9B61;
    (* HLUTNM = "LUT62_1_68" *)
    LUT2 ix12903z1488 (.O (nx12903z170), .I0 (\plaintext(54)  ), .I1 (nx34235z34
         )) ;
         defparam ix12903z1488.INIT = 4'h9;
    LUT4 ix13298z39830 (.O (nx13298z12), .I0 (\plaintext(46)  ), .I1 (
         \p_key_samp(37)  ), .I2 (nx34235z37), .I3 (nx13298z13)) ;
         defparam ix13298z39830.INIT = 16'h9669;
    LUT6 ix13298z39836 (.O (nx13298z13), .I0 (nx15291z27), .I1 (nx15291z28), .I2 (
         nx15291z30), .I3 (nx15291z31), .I4 (nx15291z33), .I5 (nx15291z34)) ;
         defparam ix13298z39836.INIT = 64'h5AA5696941B9966E;
    (* HLUTNM = "LUT62_1_67" *)
    LUT2 ix12903z1450 (.O (nx12903z134), .I0 (\plaintext(46)  ), .I1 (nx34235z37
         )) ;
         defparam ix12903z1450.INIT = 4'h6;
    (* HLUTNM = "LUT62_1_66" *)
    LUT2 ix12903z1447 (.O (nx12903z130), .I0 (\plaintext(11)  ), .I1 (nx16286z6)
         ) ;
         defparam ix12903z1447.INIT = 4'h6;
    LUT4 ix13298z28415 (.O (nx13298z71), .I0 (\plaintext(19)  ), .I1 (
         \p_key_samp(3)  ), .I2 (nx16286z9), .I3 (nx13298z72)) ;
         defparam ix13298z28415.INIT = 16'h6996;
    LUT6 ix13298z7236 (.O (nx13298z72), .I0 (nx7313z3), .I1 (nx7313z5), .I2 (
         nx7313z6), .I3 (nx7313z8), .I4 (nx7313z9), .I5 (nx7313z11)) ;
         defparam ix13298z7236.INIT = 64'h2BC7BC34D42A16DA;
    LUT4 ix7313z28354 (.O (nx7313z11), .I0 (\plaintext(34)  ), .I1 (
         \p_key_samp(11)  ), .I2 (nx41222z2), .I3 (px3688)) ;
         defparam ix7313z28354.INIT = 16'h6996;
    LUT6 ix7313z9121 (.O (px3688), .I0 (nx34235z3), .I1 (nx34235z5), .I2 (
         nx34235z7), .I3 (nx34235z9), .I4 (nx34235z20), .I5 (nx34235z30)) ;
         defparam ix7313z9121.INIT = 64'h34DDE10BE91A1E74;
    (* HLUTNM = "LUT62_1_108" *)
    LUT2 ix41222z1323 (.O (px3689), .I0 (\plaintext(34)  ), .I1 (nx41222z2)) ;
         defparam ix41222z1323.INIT = 4'h9;
    LUT4 ix7313z39827 (.O (nx7313z9), .I0 (\plaintext(50)  ), .I1 (
         \p_key_samp(51)  ), .I2 (nx34235z13), .I3 (nx7313z10)) ;
         defparam ix7313z39827.INIT = 16'h9669;
    LUT6 ix7313z38968 (.O (nx7313z10), .I0 (nx15291z17), .I1 (px3697), .I2 (
         nx15291z20), .I3 (nx15291z21), .I4 (nx15291z22), .I5 (nx15291z23)) ;
         defparam ix7313z38968.INIT = 64'hA7A978D16C9A930D;
    LUT3 ix15291z1440 (.O (nx15291z23), .I0 (\plaintext(23)  ), .I1 (
         \p_key_samp(28)  ), .I2 (nx15291z24)) ;
         defparam ix15291z1440.INIT = 8'h69;
    LUT6 ix15291z32373 (.O (nx15291z24), .I0 (nx29253z3), .I1 (nx29253z5), .I2 (
         nx29253z4), .I3 (nx29253z7), .I4 (nx29253z9), .I5 (nx29253z6)) ;
         defparam ix15291z32373.INIT = 64'h966E82711EA1793D;
    LUT3 ix15291z1484 (.O (nx15291z22), .I0 (\plaintext(7)  ), .I1 (
         \p_key_samp(37)  ), .I2 (nx34235z6)) ;
         defparam ix15291z1484.INIT = 8'h96;
    LUT3 ix15291z1483 (.O (nx15291z21), .I0 (\plaintext(31)  ), .I1 (
         \p_key_samp(39)  ), .I2 (nx28253z2)) ;
         defparam ix15291z1483.INIT = 8'h96;
    LUT3 ix15291z1482 (.O (nx15291z20), .I0 (\plaintext(57)  ), .I1 (
         \p_key_samp(13)  ), .I2 (nx34235z21)) ;
         defparam ix15291z1482.INIT = 8'h96;
    LUT3 ix15291z1435 (.O (nx15291z17), .I0 (\plaintext(15)  ), .I1 (
         \p_key_samp(54)  ), .I2 (nx15291z18)) ;
         defparam ix15291z1435.INIT = 8'h69;
    LUT6 ix15291z12686 (.O (nx15291z18), .I0 (nx34235z39), .I1 (nx34235z32), .I2 (
         nx34235z38), .I3 (nx34235z36), .I4 (nx34235z33), .I5 (nx34235z35)) ;
         defparam ix15291z12686.INIT = 64'h8146D369FEA12C5B;
    (* HLUTNM = "LUT62_1_71" *)
    LUT2 ix12903z1509 (.O (nx12903z193), .I0 (\plaintext(50)  ), .I1 (nx34235z13
         )) ;
         defparam ix12903z1509.INIT = 4'h9;
    LUT4 ix7313z39826 (.O (nx7313z8), .I0 (plaintext[6]), .I1 (\p_key_samp(44)  
         ), .I2 (nx44209z2), .I3 (px3702)) ;
         defparam ix7313z39826.INIT = 16'h9669;
    LUT6 ix16286z31417 (.O (px3702), .I0 (nx16286z3), .I1 (nx16286z4), .I2 (
         nx16286z5), .I3 (nx16286z7), .I4 (nx16286z8), .I5 (nx16286z10)) ;
         defparam ix16286z31417.INIT = 64'h2CF55928A95A7596;
    (* HLUTNM = "LUT62_1_108" *)
    LUT2 ix44209z1323 (.O (px3703), .I0 (plaintext[6]), .I1 (nx44209z2)) ;
         defparam ix44209z1323.INIT = 4'h9;
    LUT4 ix7313z28349 (.O (nx7313z6), .I0 (\plaintext(58)  ), .I1 (
         \p_key_samp(18)  ), .I2 (nx34235z18), .I3 (px3705)) ;
         defparam ix7313z28349.INIT = 16'h6996;
    LUT6 ix7313z15855 (.O (px3705), .I0 (nx15291z27), .I1 (nx15291z28), .I2 (
         nx15291z30), .I3 (nx15291z31), .I4 (nx15291z33), .I5 (nx15291z34)) ;
         defparam ix7313z15855.INIT = 64'h7899972A877838C7;
    LUT3 ix15291z1451 (.O (nx15291z34), .I0 (\p_plaintext(63)  ), .I1 (
         \p_key_samp(20)  ), .I2 (nx29253z2)) ;
         defparam ix15291z1451.INIT = 8'h69;
    LUT3 ix15291z1495 (.O (nx15291z33), .I0 (\plaintext(29)  ), .I1 (
         \p_key_samp(15)  ), .I2 (nx23267z2)) ;
         defparam ix15291z1495.INIT = 8'h96;
    LUT3 ix15291z1493 (.O (nx15291z31), .I0 (\plaintext(21)  ), .I1 (
         \p_key_samp(63)  ), .I2 (nx15291z32)) ;
         defparam ix15291z1493.INIT = 8'h96;
    LUT6 ix15291z24609 (.O (nx15291z32), .I0 (nx34235z17), .I1 (nx34235z16), .I2 (
         nx34235z12), .I3 (nx34235z14), .I4 (nx34235z19), .I5 (nx34235z11)) ;
         defparam ix15291z24609.INIT = 64'h946BAD34BC165AE1;
    LUT3 ix15291z1492 (.O (nx15291z30), .I0 (\p_plaintext(37)  ), .I1 (
         \p_key_samp(30)  ), .I2 (px3745)) ;
         defparam ix15291z1492.INIT = 8'h96;
    LUT3 ix15291z1445 (.O (nx15291z28), .I0 (\plaintext(13)  ), .I1 (
         \p_key_samp(62)  ), .I2 (nx15291z29)) ;
         defparam ix15291z1445.INIT = 8'h69;
    LUT6 ix15291z24054 (.O (nx15291z29), .I0 (nx36228z3), .I1 (nx36228z5), .I2 (
         nx36228z7), .I3 (nx36228z9), .I4 (nx36228z11), .I5 (nx36228z12)) ;
         defparam ix15291z24054.INIT = 64'h519A877C2E8758B9;
    LUT3 ix15291z1489 (.O (nx15291z27), .I0 (p_nbus_plaintext[63]), .I1 (
         \p_key_samp(53)  ), .I2 (nx63157z2)) ;
         defparam ix15291z1489.INIT = 8'h96;
    (* HLUTNM = "LUT62_1_109" *)
    LUT2 ix45207z1320 (.O (px3714), .I0 (\plaintext(58)  ), .I1 (nx34235z18)) ;
         defparam ix45207z1320.INIT = 4'h6;
    LUT4 ix7313z28348 (.O (nx7313z5), .I0 (\plaintext(26)  ), .I1 (
         \p_key_samp(57)  ), .I2 (nx45210z2), .I3 (px3716)) ;
         defparam ix7313z28348.INIT = 16'h6996;
    LUT6 ix16289z21089 (.O (px3716), .I0 (nx16289z3), .I1 (nx16289z4), .I2 (
         px3744), .I3 (nx16289z6), .I4 (nx16289z8), .I5 (nx16289z9)) ;
         defparam ix16289z21089.INIT = 64'h65A6A9D35A814D3E;
    (* HLUTNM = "LUT62_1_109" *)
    LUT2 ix45210z1323 (.O (px3717), .I0 (\plaintext(26)  ), .I1 (nx45210z2)) ;
         defparam ix45210z1323.INIT = 4'h9;
    LUT4 ix7313z28346 (.O (nx7313z3), .I0 (\plaintext(42)  ), .I1 (
         \p_key_samp(1)  ), .I2 (nx34235z15), .I3 (nx7313z4)) ;
         defparam ix7313z28346.INIT = 16'h6996;
    LUT6 ix7313z32744 (.O (nx7313z4), .I0 (nx27254z12), .I1 (nx27254z6), .I2 (
         nx27254z5), .I3 (nx27254z10), .I4 (nx27254z3), .I5 (nx27254z8)) ;
         defparam ix7313z32744.INIT = 64'h5B36843DC4397AC3;
    (* HLUTNM = "LUT62_1_70" *)
    LUT2 ix12903z1503 (.O (nx12903z190), .I0 (\plaintext(42)  ), .I1 (nx34235z15
         )) ;
         defparam ix12903z1503.INIT = 4'h6;
    (* HLUTNM = "LUT62_1_69" *)
    LUT2 ix12903z1500 (.O (nx12903z186), .I0 (\plaintext(19)  ), .I1 (nx16286z9)
         ) ;
         defparam ix12903z1500.INIT = 4'h6;
    (* HLUTNM = "LUT62_1_94" *)
    LUT3 ix61487z1466 (.O (nx61487z3), .I0 (\plaintext(22)  ), .I1 (nx63157z4), 
         .I2 (nx37234z3)) ;
         defparam ix61487z1466.INIT = 8'h96;
    (* HLUTNM = "LUT62_1_32" *)
    LUT3 ix46203z1419 (.O (px3723), .I0 (p_nbus_plaintext[63]), .I1 (nx63157z2)
         , .I2 (px3724)) ;
         defparam ix46203z1419.INIT = 8'h69;
    LUT6 ix13298z19671 (.O (px3724), .I0 (nx37234z2), .I1 (nx37234z4), .I2 (
         nx37234z6), .I3 (nx37234z9), .I4 (nx37234z5), .I5 (nx37234z8)) ;
         defparam ix13298z19671.INIT = 64'h51ACBAC3A8F34794;
    LUT4 ix37234z28351 (.O (nx37234z8), .I0 (\plaintext(38)  ), .I1 (
         \p_key_samp(22)  ), .I2 (nx63157z36), .I3 (px3726)) ;
         defparam ix37234z28351.INIT = 16'h6996;
    LUT6 ix34235z32229 (.O (px3726), .I0 (nx34235z3), .I1 (nx34235z5), .I2 (
         nx34235z7), .I3 (nx34235z9), .I4 (nx34235z20), .I5 (nx34235z30)) ;
         defparam ix34235z32229.INIT = 64'hD247952EA57978C2;
    LUT3 ix34235z1493 (.O (nx34235z30), .I0 (\plaintext(25)  ), .I1 (
         \p_key_samp(43)  ), .I2 (nx34235z31)) ;
         defparam ix34235z1493.INIT = 8'h96;
    LUT3 ix34235z1483 (.O (nx34235z20), .I0 (\plaintext(57)  ), .I1 (
         \p_key_samp(33)  ), .I2 (nx34235z21)) ;
         defparam ix34235z1483.INIT = 8'h96;
    LUT6 ix34235z39903 (.O (nx34235z21), .I0 (nx34235z22), .I1 (nx34235z23), .I2 (
         nx34235z24), .I3 (nx34235z26), .I4 (nx34235z27), .I5 (nx34235z29)) ;
         defparam ix34235z39903.INIT = 64'hD9E562923C6396A9;
    LUT3 ix34235z1472 (.O (nx34235z9), .I0 (\plaintext(33)  ), .I1 (
         \p_key_samp(11)  ), .I2 (nx34235z10)) ;
         defparam ix34235z1472.INIT = 8'h96;
    LUT3 ix34235z1425 (.O (nx34235z7), .I0 (\plaintext(41)  ), .I1 (
         \p_key_samp(44)  ), .I2 (nx34235z8)) ;
         defparam ix34235z1425.INIT = 8'h69;
    LUT6 ix34235z54991 (.O (nx34235z8), .I0 (nx37232z3), .I1 (nx37232z5), .I2 (
         nx37232z7), .I3 (nx37232z8), .I4 (nx37232z10), .I5 (nx37232z12)) ;
         defparam ix34235z54991.INIT = 64'h57896596E453D1A6;
    LUT3 ix34235z1468 (.O (nx34235z5), .I0 (\plaintext(7)  ), .I1 (
         \p_key_samp(57)  ), .I2 (nx34235z6)) ;
         defparam ix34235z1468.INIT = 8'h96;
    LUT6 ix34235z26364 (.O (nx34235z6), .I0 (nx36228z3), .I1 (nx36228z5), .I2 (
         nx36228z7), .I3 (nx36228z9), .I4 (nx36228z11), .I5 (nx36228z12)) ;
         defparam ix34235z26364.INIT = 64'h67591EE0B81E61D5;
    LUT3 ix34235z1466 (.O (nx34235z3), .I0 (\plaintext(49)  ), .I1 (
         \p_key_samp(26)  ), .I2 (nx34235z4)) ;
         defparam ix34235z1466.INIT = 8'h96;
    LUT6 ix34235z59563 (.O (nx34235z4), .I0 (nx63157z27), .I1 (nx63157z43), .I2 (
         nx63157z35), .I3 (nx63157z3), .I4 (nx63157z11), .I5 (nx63157z19)) ;
         defparam ix34235z59563.INIT = 64'hE79A54291675E386;
    (* HLUTNM = "LUT62_1_110" *)
    LUT2 ix47204z1320 (.O (px3737), .I0 (\plaintext(38)  ), .I1 (nx63157z36)) ;
         defparam ix47204z1320.INIT = 4'h6;
    LUT4 ix37234z28348 (.O (nx37234z5), .I0 (plaintext[0]), .I1 (
         \p_key_samp(53)  ), .I2 (nx63157z28), .I3 (px3739)) ;
         defparam ix37234z28348.INIT = 16'h6996;
    LUT6 ix47206z32079 (.O (px3739), .I0 (nx16289z4), .I1 (nx16289z8), .I2 (
         nx16289z3), .I3 (px3744), .I4 (nx16289z6), .I5 (nx16289z9)) ;
         defparam ix47206z32079.INIT = 64'h13C9E59E9E30782D;
    LUT3 ix16289z1426 (.O (nx16289z9), .I0 (\plaintext(53)  ), .I1 (
         \p_key_samp(61)  ), .I2 (nx16289z10)) ;
         defparam ix16289z1426.INIT = 8'h69;
    LUT6 ix16289z28578 (.O (nx16289z10), .I0 (nx39226z6), .I1 (nx39226z16), .I2 (
         nx39226z3), .I3 (nx39226z18), .I4 (nx39226z5), .I5 (nx39226z14)) ;
         defparam ix16289z28578.INIT = 64'hC92B95C366B46A78;
    LUT3 ix16289z1423 (.O (nx16289z6), .I0 (\plaintext(45)  ), .I1 (
         \p_key_samp(23)  ), .I2 (nx16289z7)) ;
         defparam ix16289z1423.INIT = 8'h69;
    LUT6 ix16289z7117 (.O (nx16289z7), .I0 (nx29253z3), .I1 (nx29253z5), .I2 (
         nx29253z4), .I3 (nx29253z7), .I4 (nx29253z9), .I5 (nx29253z6)) ;
         defparam ix16289z7117.INIT = 64'hC196B6599B6916A6;
    LUT6 ix23270z27839 (.O (px3745), .I0 (nx34235z39), .I1 (nx34235z32), .I2 (
         nx34235z38), .I3 (nx34235z36), .I4 (nx34235z33), .I5 (nx34235z35)) ;
         defparam ix23270z27839.INIT = 64'hC71E38E16992679C;
    LUT3 ix16289z1466 (.O (nx16289z3), .I0 (\plaintext(29)  ), .I1 (
         \p_key_samp(29)  ), .I2 (nx23267z2)) ;
         defparam ix16289z1466.INIT = 8'h96;
    LUT6 ix23267z30390 (.O (nx23267z2), .I0 (nx34235z22), .I1 (nx34235z23), .I2 (
         nx34235z24), .I3 (nx34235z26), .I4 (nx34235z27), .I5 (nx34235z29)) ;
         defparam ix23267z30390.INIT = 64'h966336A96CC67193;
    LUT3 ix16289z1470 (.O (nx16289z8), .I0 (\plaintext(61)  ), .I1 (
         \p_key_samp(5)  ), .I2 (nx37232z2)) ;
         defparam ix16289z1470.INIT = 8'h96;
    LUT3 ix16289z1467 (.O (nx16289z4), .I0 (plaintext[3]), .I1 (\p_key_samp(47)  
         ), .I2 (nx38222z2)) ;
         defparam ix16289z1467.INIT = 8'h96;
    (* HLUTNM = "LUT62_1_110" *)
    LUT2 ix49191z1320 (.O (px3750), .I0 (plaintext[0]), .I1 (nx63157z28)) ;
         defparam ix49191z1320.INIT = 4'h6;
    LUT4 ix37234z28352 (.O (nx37234z9), .I0 (\plaintext(30)  ), .I1 (
         \p_key_samp(55)  ), .I2 (nx63157z44), .I3 (px3752)) ;
         defparam ix37234z28352.INIT = 16'h6996;
    LUT6 ix25263z53176 (.O (px3752), .I0 (nx25263z3), .I1 (nx25263z4), .I2 (
         nx25263z5), .I3 (nx25263z7), .I4 (nx25263z9), .I5 (nx25263z10)) ;
         defparam ix25263z53176.INIT = 64'hCA393DE095CACA95;
    LUT3 ix25263z1428 (.O (nx25263z10), .I0 (plaintext[5]), .I1 (
         \p_key_samp(59)  ), .I2 (nx27254z7)) ;
         defparam ix25263z1428.INIT = 8'h69;
    LUT3 ix25263z1427 (.O (nx25263z9), .I0 (\plaintext(27)  ), .I1 (
         \p_key_samp(41)  ), .I2 (nx36228z2)) ;
         defparam ix25263z1427.INIT = 8'h69;
    LUT3 ix25263z1470 (.O (nx25263z7), .I0 (\plaintext(51)  ), .I1 (
         \p_key_samp(35)  ), .I2 (nx25263z8)) ;
         defparam ix25263z1470.INIT = 8'h96;
    LUT6 ix25263z28421 (.O (nx25263z8), .I0 (nx63157z3), .I1 (nx63157z11), .I2 (
         nx63157z19), .I3 (nx63157z27), .I4 (nx63157z35), .I5 (nx63157z43)) ;
         defparam ix25263z28421.INIT = 64'h6897354A335A69DC;
    LUT3 ix25263z1468 (.O (nx25263z5), .I0 (\plaintext(43)  ), .I1 (
         \p_key_samp(52)  ), .I2 (nx25263z6)) ;
         defparam ix25263z1468.INIT = 8'h96;
    LUT6 ix25263z16107 (.O (nx25263z6), .I0 (nx34235z23), .I1 (nx34235z22), .I2 (
         nx34235z26), .I3 (nx34235z27), .I4 (nx34235z29), .I5 (nx34235z24)) ;
         defparam ix25263z16107.INIT = 64'h3D84365BC37A39C4;
    LUT3 ix25263z1467 (.O (nx25263z4), .I0 (\plaintext(35)  ), .I1 (
         \p_key_samp(58)  ), .I2 (nx39226z2)) ;
         defparam ix25263z1467.INIT = 8'h96;
    LUT3 ix25263z1421 (.O (nx25263z3), .I0 (\plaintext(59)  ), .I1 (
         \p_key_samp(2)  ), .I2 (nx27254z4)) ;
         defparam ix25263z1421.INIT = 8'h69;
    (* HLUTNM = "LUT62_1_111" *)
    LUT2 ix50189z1320 (.O (px3761), .I0 (\plaintext(30)  ), .I1 (nx63157z44)) ;
         defparam ix50189z1320.INIT = 4'h6;
    LUT4 ix37234z28349 (.O (nx37234z6), .I0 (\plaintext(14)  ), .I1 (
         \p_key_samp(5)  ), .I2 (nx63157z12), .I3 (nx37234z7)) ;
         defparam ix37234z28349.INIT = 16'h6996;
    LUT6 ix37234z20669 (.O (nx37234z7), .I0 (nx15291z5), .I1 (nx15291z6), .I2 (
         nx15291z7), .I3 (nx15291z9), .I4 (nx15291z10), .I5 (nx15291z11)) ;
         defparam ix37234z20669.INIT = 64'hB93C3666348B4B95;
    LUT3 ix15291z1474 (.O (nx15291z11), .I0 (\plaintext(47)  ), .I1 (
         \p_key_samp(21)  ), .I2 (nx15291z12)) ;
         defparam ix15291z1474.INIT = 8'h96;
    LUT6 ix15291z8162 (.O (nx15291z12), .I0 (nx37232z3), .I1 (nx37232z5), .I2 (
         nx37232z7), .I3 (nx37232z8), .I4 (nx37232z10), .I5 (nx37232z12)) ;
         defparam ix15291z8162.INIT = 64'h3CA5C35A36691AB5;
    LUT3 ix15291z1428 (.O (nx15291z10), .I0 (\p_plaintext(63)  ), .I1 (
         \p_key_samp(4)  ), .I2 (nx29253z2)) ;
         defparam ix15291z1428.INIT = 8'h69;
    LUT6 ix29253z35726 (.O (nx29253z2), .I0 (nx29253z3), .I1 (nx29253z4), .I2 (
         nx29253z5), .I3 (nx29253z6), .I4 (nx29253z7), .I5 (nx29253z9)) ;
         defparam ix29253z35726.INIT = 64'h4D923C35AB5C866B;
    LUT3 ix15291z1472 (.O (nx15291z9), .I0 (\plaintext(31)  ), .I1 (
         \p_key_samp(55)  ), .I2 (nx28253z2)) ;
         defparam ix15291z1472.INIT = 8'h96;
    LUT6 ix28253z29004 (.O (nx28253z2), .I0 (nx34235z17), .I1 (nx34235z16), .I2 (
         nx34235z12), .I3 (nx34235z14), .I4 (nx34235z19), .I5 (nx34235z11)) ;
         defparam ix28253z29004.INIT = 64'h3D56D32DC2966C29;
    LUT3 ix15291z1425 (.O (nx15291z7), .I0 (\plaintext(55)  ), .I1 (
         \p_key_samp(14)  ), .I2 (nx15291z8)) ;
         defparam ix15291z1425.INIT = 8'h69;
    LUT6 ix15291z7411 (.O (nx15291z8), .I0 (nx34235z22), .I1 (nx34235z23), .I2 (
         nx34235z24), .I3 (nx34235z26), .I4 (nx34235z27), .I5 (nx34235z29)) ;
         defparam ix15291z7411.INIT = 64'h1EC96935C93617CA;
    LUT3 ix34235z1492 (.O (nx34235z29), .I0 (\plaintext(58)  ), .I1 (
         \p_key_samp(11)  ), .I2 (nx34235z18)) ;
         defparam ix34235z1492.INIT = 8'h96;
    LUT3 ix34235z1445 (.O (nx34235z27), .I0 (\plaintext(16)  ), .I1 (
         \p_key_samp(9)  ), .I2 (nx34235z28)) ;
         defparam ix34235z1445.INIT = 8'h69;
    LUT6 ix34235z53732 (.O (nx34235z28), .I0 (nx63157z41), .I1 (nx63157z40), .I2 (
         nx63157z37), .I3 (nx63157z38), .I4 (nx63157z42), .I5 (nx63157z39)) ;
         defparam ix34235z53732.INIT = 64'h0FE19378721CCCA7;
    LUT3 ix34235z1489 (.O (nx34235z26), .I0 (\plaintext(32)  ), .I1 (
         \p_key_samp(52)  ), .I2 (nx39226z15)) ;
         defparam ix34235z1489.INIT = 8'h96;
    LUT3 ix34235z1487 (.O (nx34235z24), .I0 (\plaintext(8)  ), .I1 (
         \p_key_samp(34)  ), .I2 (nx34235z25)) ;
         defparam ix34235z1487.INIT = 8'h96;
    LUT6 ix34235z20622 (.O (nx34235z25), .I0 (nx63157z29), .I1 (nx63157z30), .I2 (
         nx63157z31), .I3 (nx63157z32), .I4 (nx63157z33), .I5 (nx63157z34)) ;
         defparam ix34235z20622.INIT = 64'hD6B91DE2A1874B54;
    LUT3 ix34235z1441 (.O (nx34235z23), .I0 (\plaintext(24)  ), .I1 (
         \p_key_samp(57)  ), .I2 (nx39226z17)) ;
         defparam ix34235z1441.INIT = 8'h69;
    LUT3 ix34235z1440 (.O (nx34235z22), .I0 (plaintext[6]), .I1 (
         \p_key_samp(51)  ), .I2 (nx44209z2)) ;
         defparam ix34235z1440.INIT = 8'h69;
    LUT3 ix15291z1469 (.O (nx15291z6), .I0 (\p_plaintext(39)  ), .I1 (
         \p_key_samp(31)  ), .I2 (px3781)) ;
         defparam ix15291z1469.INIT = 8'h96;
    LUT6 ix28250z35919 (.O (px3781), .I0 (nx39226z3), .I1 (nx39226z5), .I2 (
         nx39226z6), .I3 (nx39226z14), .I4 (nx39226z16), .I5 (nx39226z18)) ;
         defparam ix28250z35919.INIT = 64'h2D745A9759E2872C;
    LUT3 ix15291z1468 (.O (nx15291z5), .I0 (p_nbus_plaintext[63]), .I1 (
         \p_key_samp(46)  ), .I2 (nx63157z2)) ;
         defparam ix15291z1468.INIT = 8'h96;
    (* HLUTNM = "LUT62_1_84" *)
    LUT2 ix12903z1627 (.O (nx12903z343), .I0 (\plaintext(14)  ), .I1 (nx63157z12
         )) ;
         defparam ix12903z1627.INIT = 4'h9;
    LUT4 ix37234z28347 (.O (nx37234z4), .I0 (\plaintext(56)  ), .I1 (
         \p_key_samp(29)  ), .I2 (nx63157z20), .I3 (nx27254z2)) ;
         defparam ix37234z28347.INIT = 16'h6996;
    LUT6 ix27254z49482 (.O (nx27254z2), .I0 (nx27254z3), .I1 (nx27254z5), .I2 (
         nx27254z6), .I3 (nx27254z8), .I4 (nx27254z10), .I5 (nx27254z12)) ;
         defparam ix27254z49482.INIT = 64'hB42857C969D2BC27;
    LUT3 ix27254z1475 (.O (nx27254z12), .I0 (\plaintext(25)  ), .I1 (
         \p_key_samp(10)  ), .I2 (nx34235z31)) ;
         defparam ix27254z1475.INIT = 8'h96;
    LUT6 ix34235z41460 (.O (nx34235z31), .I0 (nx34235z32), .I1 (nx34235z33), .I2 (
         nx34235z35), .I3 (nx34235z36), .I4 (nx34235z38), .I5 (nx34235z39)) ;
         defparam ix34235z41460.INIT = 64'hDC86235B23799CB4;
    LUT3 ix27254z1428 (.O (nx27254z10), .I0 (\plaintext(17)  ), .I1 (
         \p_key_samp(25)  ), .I2 (nx27254z11)) ;
         defparam ix27254z1428.INIT = 8'h69;
    LUT6 ix27254z27586 (.O (nx27254z11), .I0 (nx39226z3), .I1 (nx39226z5), .I2 (
         nx39226z6), .I3 (nx39226z14), .I4 (nx39226z16), .I5 (nx39226z18)) ;
         defparam ix27254z27586.INIT = 64'h8768C399749B6696;
    LUT3 ix27254z1471 (.O (nx27254z8), .I0 (\plaintext(9)  ), .I1 (
         \p_key_samp(50)  ), .I2 (nx27254z9)) ;
         defparam ix27254z1471.INIT = 8'h96;
    LUT6 ix27254z3234 (.O (nx27254z9), .I0 (nx36228z3), .I1 (nx36228z5), .I2 (
         nx36228z7), .I3 (nx36228z9), .I4 (nx36228z11), .I5 (nx36228z12)) ;
         defparam ix27254z3234.INIT = 64'h781DAB869AE60778;
    LUT3 ix27254z1424 (.O (nx27254z6), .I0 (plaintext[5]), .I1 (\p_key_samp(36)  
         ), .I2 (nx27254z7)) ;
         defparam ix27254z1424.INIT = 8'h69;
    LUT6 ix27254z9496 (.O (nx27254z7), .I0 (nx29253z3), .I1 (nx29253z5), .I2 (
         nx29253z4), .I3 (nx29253z7), .I4 (nx29253z9), .I5 (nx29253z6)) ;
         defparam ix27254z9496.INIT = 64'h983A61C727C91FF0;
    LUT3 ix29253z1469 (.O (nx29253z6), .I0 (plaintext[4]), .I1 (\p_key_samp(44)  
         ), .I2 (nx36228z6)) ;
         defparam ix29253z1469.INIT = 8'h96;
    LUT3 ix29253z1427 (.O (nx29253z9), .I0 (\plaintext(10)  ), .I1 (
         \p_key_samp(33)  ), .I2 (nx29253z10)) ;
         defparam ix29253z1427.INIT = 8'h69;
    LUT6 ix29253z15879 (.O (nx29253z10), .I0 (nx63157z13), .I1 (nx63157z15), .I2 (
         nx63157z18), .I3 (nx63157z16), .I4 (nx63157z14), .I5 (px3923)) ;
         defparam ix29253z15879.INIT = 64'h4AF55B286D2338DC;
    LUT3 ix29253z1470 (.O (nx29253z7), .I0 (\plaintext(18)  ), .I1 (
         \p_key_samp(18)  ), .I2 (nx29253z8)) ;
         defparam ix29253z1470.INIT = 8'h96;
    LUT6 ix29253z27278 (.O (nx29253z8), .I0 (nx63157z45), .I1 (nx63157z46), .I2 (
         nx63157z47), .I3 (nx63157z48), .I4 (nx63157z49), .I5 (nx63157z50)) ;
         defparam ix29253z27278.INIT = 64'h639CC93A8B396565;
    LUT3 ix29253z1422 (.O (nx29253z4), .I0 (\plaintext(60)  ), .I1 (
         \p_key_samp(50)  ), .I2 (nx36228z10)) ;
         defparam ix29253z1422.INIT = 8'h69;
    LUT3 ix29253z1423 (.O (nx29253z5), .I0 (\plaintext(26)  ), .I1 (
         \p_key_samp(35)  ), .I2 (nx45210z2)) ;
         defparam ix29253z1423.INIT = 8'h69;
    LUT3 ix29253z1421 (.O (nx29253z3), .I0 (\plaintext(34)  ), .I1 (
         \p_key_samp(1)  ), .I2 (nx41222z2)) ;
         defparam ix29253z1421.INIT = 8'h69;
    LUT3 ix27254z1468 (.O (nx27254z5), .I0 (\plaintext(33)  ), .I1 (
         \p_key_samp(1)  ), .I2 (nx34235z10)) ;
         defparam ix27254z1468.INIT = 8'h96;
    LUT6 ix34235z7183 (.O (nx34235z10), .I0 (nx34235z11), .I1 (nx34235z12), .I2 (
         nx34235z14), .I3 (nx34235z16), .I4 (nx34235z17), .I5 (nx34235z19)) ;
         defparam ix34235z7183.INIT = 64'h95E2E11EE95A16E4;
    LUT3 ix27254z1421 (.O (nx27254z3), .I0 (\plaintext(59)  ), .I1 (
         \p_key_samp(27)  ), .I2 (nx27254z4)) ;
         defparam ix27254z1421.INIT = 8'h69;
    LUT6 ix27254z51042 (.O (nx27254z4), .I0 (nx37232z7), .I1 (nx37232z3), .I2 (
         nx37232z10), .I3 (nx37232z5), .I4 (nx37232z12), .I5 (nx37232z8)) ;
         defparam ix27254z51042.INIT = 64'hD2662DD26D8AC23D;
    (* HLUTNM = "LUT62_1_78" *)
    LUT2 ix12903z1590 (.O (nx12903z296), .I0 (\plaintext(56)  ), .I1 (nx63157z20
         )) ;
         defparam ix12903z1590.INIT = 4'h6;
    LUT4 ix37234z28345 (.O (nx37234z2), .I0 (\plaintext(22)  ), .I1 (
         \p_key_samp(15)  ), .I2 (nx63157z4), .I3 (nx37234z3)) ;
         defparam ix37234z28345.INIT = 16'h6996;
    LUT6 ix37234z26832 (.O (nx37234z3), .I0 (nx16286z3), .I1 (nx16286z4), .I2 (
         nx16286z5), .I3 (nx16286z7), .I4 (nx16286z8), .I5 (nx16286z10)) ;
         defparam ix37234z26832.INIT = 64'hA5D9B867C60363AC;
    LUT3 ix16286z1428 (.O (nx16286z10), .I0 (\plaintext(27)  ), .I1 (
         \p_key_samp(51)  ), .I2 (nx36228z2)) ;
         defparam ix16286z1428.INIT = 8'h69;
    LUT6 ix36228z17412 (.O (nx36228z2), .I0 (nx36228z3), .I1 (nx36228z5), .I2 (
         nx36228z7), .I3 (nx36228z9), .I4 (nx36228z11), .I5 (nx36228z12)) ;
         defparam ix36228z17412.INIT = 64'hE1749D1A598A3EE1;
    LUT3 ix36228z1430 (.O (nx36228z12), .I0 (\plaintext(28)  ), .I1 (
         \p_key_samp(13)  ), .I2 (nx37232z9)) ;
         defparam ix36228z1430.INIT = 8'h69;
    LUT3 ix36228z1474 (.O (nx36228z11), .I0 (\plaintext(36)  ), .I1 (
         \p_key_samp(6)  ), .I2 (nx37232z11)) ;
         defparam ix36228z1474.INIT = 8'h96;
    LUT3 ix36228z1427 (.O (nx36228z9), .I0 (\plaintext(60)  ), .I1 (
         \p_key_samp(54)  ), .I2 (nx36228z10)) ;
         defparam ix36228z1427.INIT = 8'h69;
    LUT6 ix36228z14726 (.O (nx36228z10), .I0 (nx39226z8), .I1 (px3872), .I2 (
         nx39226z10), .I3 (px3870), .I4 (nx39226z12), .I5 (nx39226z13)) ;
         defparam ix36228z14726.INIT = 64'h16E9CB349E49345B;
    LUT3 ix36228z1425 (.O (nx36228z7), .I0 (\plaintext(52)  ), .I1 (
         \p_key_samp(45)  ), .I2 (nx36228z8)) ;
         defparam ix36228z1425.INIT = 8'h69;
    LUT6 ix36228z14517 (.O (nx36228z8), .I0 (nx63157z37), .I1 (nx63157z38), .I2 (
         nx63157z39), .I3 (nx63157z40), .I4 (nx63157z41), .I5 (nx63157z42)) ;
         defparam ix36228z14517.INIT = 64'h9625D999C679338C;
    LUT3 ix36228z1468 (.O (nx36228z5), .I0 (plaintext[4]), .I1 (\p_key_samp(31)  
         ), .I2 (nx36228z6)) ;
         defparam ix36228z1468.INIT = 8'h96;
    LUT6 ix36228z34691 (.O (nx36228z6), .I0 (nx40221z3), .I1 (nx40221z4), .I2 (
         nx40221z5), .I3 (nx40221z6), .I4 (nx40221z7), .I5 (nx40221z8)) ;
         defparam ix36228z34691.INIT = 64'h1BEC7682E769825C;
    LUT3 ix36228z1421 (.O (nx36228z3), .I0 (\plaintext(44)  ), .I1 (
         \p_key_samp(7)  ), .I2 (nx36228z4)) ;
         defparam ix36228z1421.INIT = 8'h69;
    LUT6 ix36228z35678 (.O (nx36228z4), .I0 (nx63157z7), .I1 (nx63157z5), .I2 (
         nx63157z6), .I3 (nx63157z10), .I4 (nx63157z8), .I5 (nx63157z9)) ;
         defparam ix36228z35678.INIT = 64'hA1795BC66DC28639;
    LUT3 ix16286z1471 (.O (nx16286z8), .I0 (\plaintext(19)  ), .I1 (
         \p_key_samp(34)  ), .I2 (nx16286z9)) ;
         defparam ix16286z1471.INIT = 8'h96;
    LUT6 ix16286z16022 (.O (nx16286z9), .I0 (nx34235z17), .I1 (nx34235z16), .I2 (
         nx34235z12), .I3 (nx34235z14), .I4 (nx34235z19), .I5 (nx34235z11)) ;
         defparam ix16286z16022.INIT = 64'h5A7AC5932AC5396C;
    LUT3 ix34235z1429 (.O (nx34235z11), .I0 (\plaintext(34)  ), .I1 (
         \p_key_samp(42)  ), .I2 (nx41222z2)) ;
         defparam ix34235z1429.INIT = 8'h69;
    LUT6 ix41222z24297 (.O (nx41222z2), .I0 (nx63157z37), .I1 (nx63157z38), .I2 (
         nx63157z39), .I3 (nx63157z40), .I4 (nx63157z41), .I5 (nx63157z42)) ;
         defparam ix41222z24297.INIT = 64'h1BC4E42BB23E59C6;
    LUT3 ix34235z1437 (.O (nx34235z19), .I0 (\plaintext(26)  ), .I1 (
         \p_key_samp(25)  ), .I2 (nx45210z2)) ;
         defparam ix34235z1437.INIT = 8'h69;
    LUT6 ix45210z55232 (.O (nx45210z2), .I0 (nx63157z29), .I1 (nx63157z30), .I2 (
         nx63157z31), .I3 (nx63157z32), .I4 (nx63157z33), .I5 (nx63157z34)) ;
         defparam ix45210z55232.INIT = 64'hB52A8B7468E1D29D;
    LUT3 ix34235z1477 (.O (nx34235z14), .I0 (\plaintext(42)  ), .I1 (
         \p_key_samp(36)  ), .I2 (nx34235z15)) ;
         defparam ix34235z1477.INIT = 8'h96;
    LUT6 ix34235z51561 (.O (nx34235z15), .I0 (nx63157z25), .I1 (nx63157z21), .I2 (
         nx63157z23), .I3 (nx63157z26), .I4 (nx63157z24), .I5 (nx63157z22)) ;
         defparam ix34235z51561.INIT = 64'h843D5B367AC3C439;
    LUT3 ix34235z1430 (.O (nx34235z12), .I0 (\plaintext(50)  ), .I1 (
         \p_key_samp(19)  ), .I2 (nx34235z13)) ;
         defparam ix34235z1430.INIT = 8'h69;
    LUT6 ix34235z21172 (.O (nx34235z13), .I0 (nx40221z5), .I1 (nx40221z8), .I2 (
         nx40221z4), .I3 (nx40221z3), .I4 (nx40221z6), .I5 (nx40221z7)) ;
         defparam ix34235z21172.INIT = 64'hE35AB83C17694D86;
    LUT3 ix34235z1434 (.O (nx34235z16), .I0 (plaintext[6]), .I1 (
         \p_key_samp(43)  ), .I2 (nx44209z2)) ;
         defparam ix34235z1434.INIT = 8'h69;
    LUT6 ix44209z43839 (.O (nx44209z2), .I0 (nx63157z5), .I1 (nx63157z6), .I2 (
         nx63157z7), .I3 (nx63157z8), .I4 (nx63157z9), .I5 (nx63157z10)) ;
         defparam ix44209z43839.INIT = 64'h6966D2D13C9DA61C;
    LUT3 ix34235z1480 (.O (nx34235z17), .I0 (\plaintext(58)  ), .I1 (
         \p_key_samp(49)  ), .I2 (nx34235z18)) ;
         defparam ix34235z1480.INIT = 8'h96;
    LUT6 ix34235z57192 (.O (nx34235z18), .I0 (nx39226z10), .I1 (px3872), .I2 (
         nx39226z8), .I3 (nx39226z12), .I4 (nx39226z13), .I5 (px3870)) ;
         defparam ix34235z57192.INIT = 64'h87693CC3689ADA35;
    LUT3 ix16286z1470 (.O (nx16286z7), .I0 (\plaintext(61)  ), .I1 (
         \p_key_samp(3)  ), .I2 (nx37232z2)) ;
         defparam ix16286z1470.INIT = 8'h96;
    LUT6 ix37232z23470 (.O (nx37232z2), .I0 (nx37232z3), .I1 (nx37232z5), .I2 (
         nx37232z7), .I3 (nx37232z8), .I4 (nx37232z10), .I5 (nx37232z12)) ;
         defparam ix37232z23470.INIT = 64'h7A43297CA53C568B;
    LUT3 ix37232z1475 (.O (nx37232z12), .I0 (\plaintext(62)  ), .I1 (
         \p_key_samp(4)  ), .I2 (nx37232z13)) ;
         defparam ix37232z1475.INIT = 8'h96;
    LUT3 ix37232z1473 (.O (nx37232z10), .I0 (\plaintext(36)  ), .I1 (
         \p_key_samp(14)  ), .I2 (nx37232z11)) ;
         defparam ix37232z1473.INIT = 8'h96;
    LUT6 ix37232z39806 (.O (nx37232z11), .I0 (nx63157z13), .I1 (nx63157z14), .I2 (
         nx63157z15), .I3 (nx63157z16), .I4 (px3923), .I5 (nx63157z18)) ;
         defparam ix37232z39806.INIT = 64'h39D266AD668D9652;
    LUT3 ix37232z1426 (.O (nx37232z8), .I0 (\plaintext(28)  ), .I1 (
         \p_key_samp(28)  ), .I2 (nx37232z9)) ;
         defparam ix37232z1426.INIT = 8'h69;
    LUT6 ix37232z39335 (.O (nx37232z9), .I0 (nx63157z21), .I1 (nx63157z22), .I2 (
         nx63157z23), .I3 (nx63157z24), .I4 (nx63157z25), .I5 (nx63157z26)) ;
         defparam ix37232z39335.INIT = 64'hE5B716286B82947D;
    LUT3 ix37232z1470 (.O (nx37232z7), .I0 (plaintext[2]), .I1 (\p_key_samp(37)  
         ), .I2 (nx40221z2)) ;
         defparam ix37232z1470.INIT = 8'h96;
    LUT3 ix37232z1468 (.O (nx37232z5), .I0 (\plaintext(20)  ), .I1 (
         \p_key_samp(47)  ), .I2 (nx37232z6)) ;
         defparam ix37232z1468.INIT = 8'h96;
    LUT6 ix37232z40199 (.O (nx37232z6), .I0 (nx63157z45), .I1 (nx63157z46), .I2 (
         nx63157z47), .I3 (nx63157z48), .I4 (nx63157z49), .I5 (nx63157z50)) ;
         defparam ix37232z40199.INIT = 64'h39E94E164A9797E0;
    LUT3 ix37232z1466 (.O (nx37232z3), .I0 (\plaintext(12)  ), .I1 (
         \p_key_samp(46)  ), .I2 (nx37232z4)) ;
         defparam ix37232z1466.INIT = 8'h96;
    LUT6 ix37232z44419 (.O (nx37232z4), .I0 (nx63157z29), .I1 (nx63157z30), .I2 (
         nx63157z31), .I3 (nx63157z32), .I4 (nx63157z33), .I5 (nx63157z34)) ;
         defparam ix37232z44419.INIT = 64'h76874B291DE2A85E;
    LUT3 ix16286z1468 (.O (nx16286z5), .I0 (\plaintext(11)  ), .I1 (
         \p_key_samp(49)  ), .I2 (nx16286z6)) ;
         defparam ix16286z1468.INIT = 8'h96;
    LUT6 ix16286z54281 (.O (nx16286z6), .I0 (nx34235z39), .I1 (nx34235z32), .I2 (
         nx34235z38), .I3 (nx34235z36), .I4 (nx34235z33), .I5 (nx34235z35)) ;
         defparam ix16286z54281.INIT = 64'hE28D523D3915CEE2;
    LUT3 ix34235z1498 (.O (nx34235z35), .I0 (\plaintext(38)  ), .I1 (
         \p_key_samp(15)  ), .I2 (nx63157z36)) ;
         defparam ix34235z1498.INIT = 8'h96;
    LUT3 ix34235z1451 (.O (nx34235z33), .I0 (\plaintext(54)  ), .I1 (
         \p_key_samp(63)  ), .I2 (nx34235z34)) ;
         defparam ix34235z1451.INIT = 8'h69;
    LUT6 ix34235z58977 (.O (nx34235z34), .I0 (nx63157z21), .I1 (nx63157z22), .I2 (
         nx63157z25), .I3 (nx63157z23), .I4 (nx63157z26), .I5 (nx63157z24)) ;
         defparam ix34235z58977.INIT = 64'h691D36E117E2E11E;
    LUT3 ix34235z1499 (.O (nx34235z36), .I0 (\plaintext(46)  ), .I1 (
         \p_key_samp(5)  ), .I2 (nx34235z37)) ;
         defparam ix34235z1499.INIT = 8'h96;
    LUT6 ix34235z8924 (.O (nx34235z37), .I0 (nx39226z8), .I1 (px3872), .I2 (
         nx39226z10), .I3 (px3870), .I4 (nx39226z12), .I5 (nx39226z13)) ;
         defparam ix34235z8924.INIT = 64'h6DC35296D23C1D96;
    LUT3 ix34235z1501 (.O (nx34235z38), .I0 (\plaintext(62)  ), .I1 (
         \p_key_samp(53)  ), .I2 (nx37232z13)) ;
         defparam ix34235z1501.INIT = 8'h96;
    LUT6 ix37232z9089 (.O (nx37232z13), .I0 (nx63157z5), .I1 (nx63157z6), .I2 (
         nx63157z7), .I3 (nx63157z8), .I4 (nx63157z9), .I5 (nx63157z10)) ;
         defparam ix37232z9089.INIT = 64'h9849E6B9A63C1E53;
    LUT3 ix34235z1495 (.O (nx34235z32), .I0 (plaintext[2]), .I1 (
         \p_key_samp(30)  ), .I2 (nx40221z2)) ;
         defparam ix34235z1495.INIT = 8'h96;
    LUT6 ix40221z52876 (.O (nx40221z2), .I0 (nx40221z3), .I1 (nx40221z4), .I2 (
         nx40221z5), .I3 (nx40221z6), .I4 (nx40221z7), .I5 (nx40221z8)) ;
         defparam ix40221z52876.INIT = 64'h826997BC935AC969;
    LUT3 ix34235z1502 (.O (nx34235z39), .I0 (\plaintext(30)  ), .I1 (
         \p_key_samp(39)  ), .I2 (nx63157z44)) ;
         defparam ix34235z1502.INIT = 8'h96;
    LUT3 ix16286z1467 (.O (nx16286z4), .I0 (\plaintext(35)  ), .I1 (
         \p_key_samp(17)  ), .I2 (nx39226z2)) ;
         defparam ix16286z1467.INIT = 8'h96;
    LUT6 ix39226z9179 (.O (nx39226z2), .I0 (nx39226z3), .I1 (nx39226z5), .I2 (
         nx39226z6), .I3 (nx39226z14), .I4 (nx39226z16), .I5 (nx39226z18)) ;
         defparam ix39226z9179.INIT = 64'hBC22615EE14F1EB8;
    LUT3 ix39226z1479 (.O (nx39226z18), .I0 (\plaintext(56)  ), .I1 (
         \p_key_samp(17)  ), .I2 (nx63157z20)) ;
         defparam ix39226z1479.INIT = 8'h96;
    LUT3 ix39226z1432 (.O (nx39226z16), .I0 (\plaintext(24)  ), .I1 (
         \p_key_samp(27)  ), .I2 (nx39226z17)) ;
         defparam ix39226z1432.INIT = 8'h69;
    LUT6 ix39226z10950 (.O (nx39226z17), .I0 (nx63157z13), .I1 (nx63157z14), .I2 (
         nx63157z15), .I3 (nx63157z16), .I4 (px3923), .I5 (nx63157z18)) ;
         defparam ix39226z10950.INIT = 64'h96967A961EE12596;
    LUT3 ix39226z1475 (.O (nx39226z14), .I0 (\plaintext(32)  ), .I1 (
         \p_key_samp(58)  ), .I2 (nx39226z15)) ;
         defparam ix39226z1475.INIT = 8'h96;
    LUT6 ix39226z43927 (.O (nx39226z15), .I0 (nx63157z49), .I1 (nx63157z48), .I2 (
         nx63157z50), .I3 (nx63157z47), .I4 (nx63157z46), .I5 (nx63157z45)) ;
         defparam ix39226z43927.INIT = 64'hB1CB4CB6433CA669;
    LUT3 ix39226z1469 (.O (nx39226z6), .I0 (\plaintext(40)  ), .I1 (
         \p_key_samp(59)  ), .I2 (nx39226z7)) ;
         defparam ix39226z1469.INIT = 8'h96;
    LUT6 ix39226z46441 (.O (nx39226z7), .I0 (nx39226z8), .I1 (px3872), .I2 (
         nx39226z10), .I3 (px3870), .I4 (nx39226z12), .I5 (nx39226z13)) ;
         defparam ix39226z46441.INIT = 64'h3949E6BFC5A6B041;
    LUT2 ix39226z1330 (.O (nx39226z13), .I0 (\plaintext(13)  ), .I1 (
         \p_key_samp(38)  )) ;
         defparam ix39226z1330.INIT = 4'h6;
    LUT2 ix39226z1329 (.O (nx39226z12), .I0 (\plaintext(29)  ), .I1 (
         \p_key_samp(20)  )) ;
         defparam ix39226z1329.INIT = 4'h6;
    LUT2 ix39226z1328 (.O (nx39226z10), .I0 (p_nbus_plaintext[63]), .I1 (
         \p_key_samp(29)  )) ;
         defparam ix39226z1328.INIT = 4'h6;
    LUT2 ix39226z1327 (.O (nx39226z8), .I0 (\plaintext(21)  ), .I1 (
         \p_key_samp(39)  )) ;
         defparam ix39226z1327.INIT = 4'h6;
    LUT3 ix39226z1468 (.O (nx39226z5), .I0 (plaintext[0]), .I1 (\p_key_samp(41)  
         ), .I2 (nx63157z28)) ;
         defparam ix39226z1468.INIT = 8'h96;
    LUT3 ix39226z1466 (.O (nx39226z3), .I0 (\plaintext(48)  ), .I1 (
         \p_key_samp(10)  ), .I2 (nx39226z4)) ;
         defparam ix39226z1466.INIT = 8'h96;
    LUT6 ix39226z29184 (.O (nx39226z4), .I0 (nx40221z3), .I1 (nx40221z4), .I2 (
         nx40221z5), .I3 (nx40221z6), .I4 (nx40221z7), .I5 (nx40221z8)) ;
         defparam ix39226z29184.INIT = 64'h49DAB32986316CDB;
    LUT2 ix40221z1327 (.O (nx40221z8), .I0 (\plaintext(57)  ), .I1 (
         \p_key_samp(54)  )) ;
         defparam ix40221z1327.INIT = 4'h6;
    LUT2 ix40221z1326 (.O (nx40221z7), .I0 (\plaintext(15)  ), .I1 (
         \p_key_samp(30)  )) ;
         defparam ix40221z1326.INIT = 4'h6;
    LUT2 ix40221z1325 (.O (nx40221z6), .I0 (\plaintext(23)  ), .I1 (
         \p_key_samp(4)  )) ;
         defparam ix40221z1325.INIT = 4'h6;
    LUT2 ix40221z1324 (.O (nx40221z5), .I0 (\p_plaintext(39)  ), .I1 (
         \p_key_samp(47)  )) ;
         defparam ix40221z1324.INIT = 4'h6;
    LUT2 ix40221z1323 (.O (nx40221z4), .I0 (\plaintext(7)  ), .I1 (
         \p_key_samp(13)  )) ;
         defparam ix40221z1323.INIT = 4'h6;
    LUT2 ix40221z1322 (.O (nx40221z3), .I0 (\plaintext(31)  ), .I1 (
         \p_key_samp(15)  )) ;
         defparam ix40221z1322.INIT = 4'h6;
    LUT3 ix16286z1466 (.O (nx16286z3), .I0 (plaintext[3]), .I1 (\p_key_samp(60)  
         ), .I2 (nx38222z2)) ;
         defparam ix16286z1466.INIT = 8'h96;
    LUT6 ix38222z59480 (.O (nx38222z2), .I0 (nx63157z35), .I1 (nx63157z27), .I2 (
         nx63157z43), .I3 (nx63157z11), .I4 (nx63157z3), .I5 (nx63157z19)) ;
         defparam ix38222z59480.INIT = 64'hE49609DB09CEE335;
    (* HLUTNM = "LUT62_1_83" *)
    LUT2 ix12903z1622 (.O (nx12903z341), .I0 (\plaintext(22)  ), .I1 (nx63157z4)
         ) ;
         defparam ix12903z1622.INIT = 4'h6;
    (* HLUTNM = "LUT62_1_111" *)
    LUT2 ix63157z1320 (.O (px3886), .I0 (p_nbus_plaintext[63]), .I1 (nx63157z2)
         ) ;
         defparam ix63157z1320.INIT = 4'h6;
    LUT6 ix63157z61272 (.O (nx63157z2), .I0 (nx63157z3), .I1 (nx63157z11), .I2 (
         nx63157z19), .I3 (nx63157z27), .I4 (nx63157z35), .I5 (nx63157z43)) ;
         defparam ix63157z61272.INIT = 64'hE23C0CD65D8AEA35;
    LUT3 ix63157z1505 (.O (nx63157z43), .I0 (\plaintext(30)  ), .I1 (
         \p_key_samp(23)  ), .I2 (nx63157z44)) ;
         defparam ix63157z1505.INIT = 8'h96;
    LUT6 ix63157z25074 (.O (nx63157z44), .I0 (nx63157z45), .I1 (nx63157z46), .I2 (
         nx63157z47), .I3 (nx63157z48), .I4 (nx63157z49), .I5 (nx63157z50)) ;
         defparam ix63157z25074.INIT = 64'h0DA6E35C635C5CA6;
    LUT2 ix63157z1368 (.O (nx63157z50), .I0 (\plaintext(27)  ), .I1 (
         \p_key_samp(17)  )) ;
         defparam ix63157z1368.INIT = 4'h6;
    LUT2 ix63157z1367 (.O (nx63157z49), .I0 (\plaintext(51)  ), .I1 (
         \p_key_samp(11)  )) ;
         defparam ix63157z1367.INIT = 4'h6;
    LUT2 ix63157z1366 (.O (nx63157z48), .I0 (plaintext[5]), .I1 (
         \p_key_samp(35)  )) ;
         defparam ix63157z1366.INIT = 4'h6;
    LUT2 ix63157z1365 (.O (nx63157z47), .I0 (\plaintext(43)  ), .I1 (
         \p_key_samp(59)  )) ;
         defparam ix63157z1365.INIT = 4'h6;
    LUT2 ix63157z1364 (.O (nx63157z46), .I0 (\plaintext(35)  ), .I1 (
         \p_key_samp(34)  )) ;
         defparam ix63157z1364.INIT = 4'h6;
    LUT2 ix63157z1363 (.O (nx63157z45), .I0 (\plaintext(59)  ), .I1 (
         \p_key_samp(41)  )) ;
         defparam ix63157z1363.INIT = 4'h6;
    LUT3 ix63157z1497 (.O (nx63157z35), .I0 (\plaintext(38)  ), .I1 (
         \p_key_samp(55)  ), .I2 (nx63157z36)) ;
         defparam ix63157z1497.INIT = 8'h96;
    LUT6 ix63157z40875 (.O (nx63157z36), .I0 (nx63157z37), .I1 (nx63157z38), .I2 (
         nx63157z39), .I3 (nx63157z40), .I4 (nx63157z41), .I5 (nx63157z42)) ;
         defparam ix63157z40875.INIT = 64'hB94941BC27E89A67;
    LUT2 ix63157z1360 (.O (nx63157z42), .I0 (\plaintext(57)  ), .I1 (
         \p_key_samp(9)  )) ;
         defparam ix63157z1360.INIT = 4'h6;
    LUT2 ix63157z1359 (.O (nx63157z41), .I0 (\plaintext(25)  ), .I1 (
         \p_key_samp(19)  )) ;
         defparam ix63157z1359.INIT = 4'h6;
    LUT2 ix63157z1358 (.O (nx63157z40), .I0 (\plaintext(41)  ), .I1 (
         \p_key_samp(51)  )) ;
         defparam ix63157z1358.INIT = 4'h6;
    LUT2 ix63157z1357 (.O (nx63157z39), .I0 (\plaintext(7)  ), .I1 (
         \p_key_samp(33)  )) ;
         defparam ix63157z1357.INIT = 4'h6;
    LUT2 ix63157z1356 (.O (nx63157z38), .I0 (\plaintext(33)  ), .I1 (
         \p_key_samp(50)  )) ;
         defparam ix63157z1356.INIT = 4'h6;
    LUT2 ix63157z1355 (.O (nx63157z37), .I0 (\plaintext(49)  ), .I1 (
         \p_key_samp(2)  )) ;
         defparam ix63157z1355.INIT = 4'h6;
    LUT3 ix63157z1489 (.O (nx63157z27), .I0 (plaintext[0]), .I1 (
         \p_key_samp(21)  ), .I2 (nx63157z28)) ;
         defparam ix63157z1489.INIT = 8'h96;
    LUT6 ix63157z29651 (.O (nx63157z28), .I0 (nx63157z29), .I1 (nx63157z30), .I2 (
         nx63157z31), .I3 (nx63157z32), .I4 (nx63157z33), .I5 (nx63157z34)) ;
         defparam ix63157z29651.INIT = 64'h15E1D24A8B746E97;
    LUT2 ix63157z1352 (.O (nx63157z34), .I0 (\plaintext(45)  ), .I1 (
         \p_key_samp(28)  )) ;
         defparam ix63157z1352.INIT = 4'h6;
    LUT2 ix63157z1351 (.O (nx63157z33), .I0 (\plaintext(53)  ), .I1 (
         \p_key_samp(37)  )) ;
         defparam ix63157z1351.INIT = 4'h6;
    LUT2 ix63157z1350 (.O (nx63157z32), .I0 (\plaintext(29)  ), .I1 (
         \p_key_samp(5)  )) ;
         defparam ix63157z1350.INIT = 4'h6;
    LUT2 ix63157z1349 (.O (nx63157z31), .I0 (\plaintext(61)  ), .I1 (
         \p_key_samp(46)  )) ;
         defparam ix63157z1349.INIT = 4'h6;
    LUT2 ix63157z1348 (.O (nx63157z30), .I0 (plaintext[3]), .I1 (
         \p_key_samp(23)  )) ;
         defparam ix63157z1348.INIT = 4'h6;
    LUT2 ix63157z1347 (.O (nx63157z29), .I0 (\p_plaintext(37)  ), .I1 (
         \p_key_samp(63)  )) ;
         defparam ix63157z1347.INIT = 4'h6;
    LUT3 ix63157z1481 (.O (nx63157z19), .I0 (\plaintext(56)  ), .I1 (
         \p_key_samp(62)  ), .I2 (nx63157z20)) ;
         defparam ix63157z1481.INIT = 8'h96;
    LUT6 ix63157z24319 (.O (nx63157z20), .I0 (nx63157z21), .I1 (nx63157z22), .I2 (
         nx63157z23), .I3 (nx63157z24), .I4 (nx63157z25), .I5 (nx63157z26)) ;
         defparam ix63157z24319.INIT = 64'h489AA669ED3459CB;
    LUT2 ix63157z1344 (.O (nx63157z26), .I0 (\plaintext(17)  ), .I1 (
         \p_key_samp(1)  )) ;
         defparam ix63157z1344.INIT = 4'h6;
    LUT2 ix63157z1343 (.O (nx63157z25), .I0 (\plaintext(25)  ), .I1 (
         \p_key_samp(49)  )) ;
         defparam ix63157z1343.INIT = 4'h6;
    LUT2 ix63157z1342 (.O (nx63157z24), .I0 (\plaintext(59)  ), .I1 (
         \p_key_samp(3)  )) ;
         defparam ix63157z1342.INIT = 4'h6;
    LUT2 ix63157z1341 (.O (nx63157z23), .I0 (\plaintext(33)  ), .I1 (
         \p_key_samp(44)  )) ;
         defparam ix63157z1341.INIT = 4'h6;
    LUT2 ix63157z1340 (.O (nx63157z22), .I0 (\plaintext(9)  ), .I1 (
         \p_key_samp(26)  )) ;
         defparam ix63157z1340.INIT = 4'h6;
    LUT2 ix63157z1339 (.O (nx63157z21), .I0 (plaintext[5]), .I1 (
         \p_key_samp(43)  )) ;
         defparam ix63157z1339.INIT = 4'h6;
    LUT3 ix63157z1429 (.O (nx63157z11), .I0 (\plaintext(14)  ), .I1 (
         \p_key_samp(38)  ), .I2 (nx63157z12)) ;
         defparam ix63157z1429.INIT = 8'h69;
    LUT6 ix63157z35862 (.O (nx63157z12), .I0 (nx63157z13), .I1 (nx63157z14), .I2 (
         nx63157z15), .I3 (nx63157z16), .I4 (px3923), .I5 (nx63157z18)) ;
         defparam ix63157z35862.INIT = 64'h45BBE817784986E9;
    LUT2 ix63157z1336 (.O (nx63157z18), .I0 (\plaintext(47)  ), .I1 (
         \p_key_samp(62)  )) ;
         defparam ix63157z1336.INIT = 4'h6;
    LUT2 ix63157z1335 (.O (nx63157z16), .I0 (\p_plaintext(39)  ), .I1 (
         \p_key_samp(7)  )) ;
         defparam ix63157z1335.INIT = 4'h6;
    LUT2 ix63157z1334 (.O (nx63157z15), .I0 (\plaintext(31)  ), .I1 (
         \p_key_samp(31)  )) ;
         defparam ix63157z1334.INIT = 4'h6;
    LUT2 ix63157z1333 (.O (nx63157z14), .I0 (\plaintext(55)  ), .I1 (
         \p_key_samp(55)  )) ;
         defparam ix63157z1333.INIT = 4'h6;
    LUT2 ix63157z1332 (.O (nx63157z13), .I0 (\p_plaintext(63)  ), .I1 (
         \p_key_samp(45)  )) ;
         defparam ix63157z1332.INIT = 4'h6;
    LUT3 ix63157z1466 (.O (nx63157z3), .I0 (\plaintext(22)  ), .I1 (
         \p_key_samp(12)  ), .I2 (nx63157z4)) ;
         defparam ix63157z1466.INIT = 8'h96;
    LUT6 ix63157z39098 (.O (nx63157z4), .I0 (nx63157z5), .I1 (nx63157z6), .I2 (
         nx63157z7), .I3 (nx63157z8), .I4 (nx63157z9), .I5 (nx63157z10)) ;
         defparam ix63157z39098.INIT = 64'h0BA17CCBD42B9395;
    LUT2 ix63157z1329 (.O (nx63157z10), .I0 (\plaintext(61)  ), .I1 (
         \p_key_samp(42)  )) ;
         defparam ix63157z1329.INIT = 4'h6;
    LUT2 ix63157z1328 (.O (nx63157z9), .I0 (\plaintext(27)  ), .I1 (
         \p_key_samp(27)  )) ;
         defparam ix63157z1328.INIT = 4'h6;
    LUT2 ix63157z1327 (.O (nx63157z8), .I0 (\plaintext(35)  ), .I1 (
         \p_key_samp(60)  )) ;
         defparam ix63157z1327.INIT = 4'h6;
    LUT2 ix63157z1326 (.O (nx63157z7), .I0 (\plaintext(19)  ), .I1 (
         \p_key_samp(10)  )) ;
         defparam ix63157z1326.INIT = 4'h6;
    LUT2 ix63157z1325 (.O (nx63157z6), .I0 (plaintext[3]), .I1 (\p_key_samp(36)  
         )) ;
         defparam ix63157z1325.INIT = 4'h6;
    LUT2 ix63157z1324 (.O (nx63157z5), .I0 (\plaintext(11)  ), .I1 (
         \p_key_samp(25)  )) ;
         defparam ix63157z1324.INIT = 4'h6;
endmodule

